
module register ( clk, rst_n, RegWrite, ReadReg1, ReadReg2, WriteReg, 
        WriteData, ReadData1, ReadData2 );
  input [4:0] ReadReg1;
  input [4:0] ReadReg2;
  input [4:0] WriteReg;
  input [31:0] WriteData;
  output [31:0] ReadData1;
  output [31:0] ReadData2;
  input clk, rst_n, RegWrite;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, \register[31][31] ,
         \register[31][30] , \register[31][29] , \register[31][28] ,
         \register[31][27] , \register[31][26] , \register[31][25] ,
         \register[31][24] , \register[31][23] , \register[31][22] ,
         \register[31][21] , \register[31][20] , \register[31][19] ,
         \register[31][18] , \register[31][17] , \register[31][16] ,
         \register[31][15] , \register[31][14] , \register[31][13] ,
         \register[31][12] , \register[31][11] , \register[31][10] ,
         \register[31][9] , \register[31][8] , \register[31][7] ,
         \register[31][6] , \register[31][5] , \register[31][4] ,
         \register[31][3] , \register[31][2] , \register[31][1] ,
         \register[31][0] , \register[30][31] , \register[30][30] ,
         \register[30][29] , \register[30][28] , \register[30][27] ,
         \register[30][26] , \register[30][25] , \register[30][24] ,
         \register[30][23] , \register[30][22] , \register[30][21] ,
         \register[30][20] , \register[30][19] , \register[30][18] ,
         \register[30][17] , \register[30][16] , \register[30][15] ,
         \register[30][14] , \register[30][13] , \register[30][12] ,
         \register[30][11] , \register[30][10] , \register[30][9] ,
         \register[30][8] , \register[30][7] , \register[30][6] ,
         \register[30][5] , \register[30][4] , \register[30][3] ,
         \register[30][2] , \register[30][1] , \register[30][0] ,
         \register[29][31] , \register[29][30] , \register[29][29] ,
         \register[29][28] , \register[29][27] , \register[29][26] ,
         \register[29][25] , \register[29][24] , \register[29][23] ,
         \register[29][22] , \register[29][21] , \register[29][20] ,
         \register[29][19] , \register[29][18] , \register[29][17] ,
         \register[29][16] , \register[29][15] , \register[29][14] ,
         \register[29][13] , \register[29][12] , \register[29][11] ,
         \register[29][10] , \register[29][9] , \register[29][8] ,
         \register[29][7] , \register[29][6] , \register[29][5] ,
         \register[29][4] , \register[29][3] , \register[29][2] ,
         \register[29][1] , \register[29][0] , \register[28][31] ,
         \register[28][30] , \register[28][29] , \register[28][28] ,
         \register[28][27] , \register[28][26] , \register[28][25] ,
         \register[28][24] , \register[28][23] , \register[28][22] ,
         \register[28][21] , \register[28][20] , \register[28][19] ,
         \register[28][18] , \register[28][17] , \register[28][16] ,
         \register[28][15] , \register[28][14] , \register[28][13] ,
         \register[28][12] , \register[28][11] , \register[28][10] ,
         \register[28][9] , \register[28][8] , \register[28][7] ,
         \register[28][6] , \register[28][5] , \register[28][4] ,
         \register[28][3] , \register[28][2] , \register[28][1] ,
         \register[28][0] , \register[27][31] , \register[27][30] ,
         \register[27][29] , \register[27][28] , \register[27][27] ,
         \register[27][26] , \register[27][25] , \register[27][24] ,
         \register[27][23] , \register[27][22] , \register[27][21] ,
         \register[27][20] , \register[27][19] , \register[27][18] ,
         \register[27][17] , \register[27][16] , \register[27][15] ,
         \register[27][14] , \register[27][13] , \register[27][12] ,
         \register[27][11] , \register[27][10] , \register[27][9] ,
         \register[27][8] , \register[27][7] , \register[27][6] ,
         \register[27][5] , \register[27][4] , \register[27][3] ,
         \register[27][2] , \register[27][1] , \register[27][0] ,
         \register[26][31] , \register[26][30] , \register[26][29] ,
         \register[26][28] , \register[26][27] , \register[26][26] ,
         \register[26][25] , \register[26][24] , \register[26][23] ,
         \register[26][22] , \register[26][21] , \register[26][20] ,
         \register[26][19] , \register[26][18] , \register[26][17] ,
         \register[26][16] , \register[26][15] , \register[26][14] ,
         \register[26][13] , \register[26][12] , \register[26][11] ,
         \register[26][10] , \register[26][9] , \register[26][8] ,
         \register[26][7] , \register[26][6] , \register[26][5] ,
         \register[26][4] , \register[26][3] , \register[26][2] ,
         \register[26][1] , \register[26][0] , \register[25][31] ,
         \register[25][30] , \register[25][29] , \register[25][28] ,
         \register[25][27] , \register[25][26] , \register[25][25] ,
         \register[25][24] , \register[25][23] , \register[25][22] ,
         \register[25][21] , \register[25][20] , \register[25][19] ,
         \register[25][18] , \register[25][17] , \register[25][16] ,
         \register[25][15] , \register[25][14] , \register[25][13] ,
         \register[25][12] , \register[25][11] , \register[25][10] ,
         \register[25][9] , \register[25][8] , \register[25][7] ,
         \register[25][6] , \register[25][5] , \register[25][4] ,
         \register[25][3] , \register[25][2] , \register[25][1] ,
         \register[25][0] , \register[24][31] , \register[24][30] ,
         \register[24][29] , \register[24][28] , \register[24][27] ,
         \register[24][26] , \register[24][25] , \register[24][24] ,
         \register[24][23] , \register[24][22] , \register[24][21] ,
         \register[24][20] , \register[24][19] , \register[24][18] ,
         \register[24][17] , \register[24][16] , \register[24][15] ,
         \register[24][14] , \register[24][13] , \register[24][12] ,
         \register[24][11] , \register[24][10] , \register[24][9] ,
         \register[24][8] , \register[24][7] , \register[24][6] ,
         \register[24][5] , \register[24][4] , \register[24][3] ,
         \register[24][2] , \register[24][1] , \register[24][0] ,
         \register[23][31] , \register[23][30] , \register[23][29] ,
         \register[23][28] , \register[23][27] , \register[23][26] ,
         \register[23][25] , \register[23][24] , \register[23][23] ,
         \register[23][22] , \register[23][21] , \register[23][20] ,
         \register[23][19] , \register[23][18] , \register[23][17] ,
         \register[23][16] , \register[23][15] , \register[23][14] ,
         \register[23][13] , \register[23][12] , \register[23][11] ,
         \register[23][10] , \register[23][9] , \register[23][8] ,
         \register[23][7] , \register[23][6] , \register[23][5] ,
         \register[23][4] , \register[23][3] , \register[23][2] ,
         \register[23][1] , \register[23][0] , \register[22][31] ,
         \register[22][30] , \register[22][29] , \register[22][28] ,
         \register[22][27] , \register[22][26] , \register[22][25] ,
         \register[22][24] , \register[22][23] , \register[22][22] ,
         \register[22][21] , \register[22][20] , \register[22][19] ,
         \register[22][18] , \register[22][17] , \register[22][16] ,
         \register[22][15] , \register[22][14] , \register[22][13] ,
         \register[22][12] , \register[22][11] , \register[22][10] ,
         \register[22][9] , \register[22][8] , \register[22][7] ,
         \register[22][6] , \register[22][5] , \register[22][4] ,
         \register[22][3] , \register[22][2] , \register[22][1] ,
         \register[22][0] , \register[21][31] , \register[21][30] ,
         \register[21][29] , \register[21][28] , \register[21][27] ,
         \register[21][26] , \register[21][25] , \register[21][24] ,
         \register[21][23] , \register[21][22] , \register[21][21] ,
         \register[21][20] , \register[21][19] , \register[21][18] ,
         \register[21][17] , \register[21][16] , \register[21][15] ,
         \register[21][14] , \register[21][13] , \register[21][12] ,
         \register[21][11] , \register[21][10] , \register[21][9] ,
         \register[21][8] , \register[21][7] , \register[21][6] ,
         \register[21][5] , \register[21][4] , \register[21][3] ,
         \register[21][2] , \register[21][1] , \register[21][0] ,
         \register[20][31] , \register[20][30] , \register[20][29] ,
         \register[20][28] , \register[20][27] , \register[20][26] ,
         \register[20][25] , \register[20][24] , \register[20][23] ,
         \register[20][22] , \register[20][21] , \register[20][20] ,
         \register[20][19] , \register[20][18] , \register[20][17] ,
         \register[20][16] , \register[20][15] , \register[20][14] ,
         \register[20][13] , \register[20][12] , \register[20][11] ,
         \register[20][10] , \register[20][9] , \register[20][8] ,
         \register[20][7] , \register[20][6] , \register[20][5] ,
         \register[20][4] , \register[20][3] , \register[20][2] ,
         \register[20][1] , \register[20][0] , \register[19][31] ,
         \register[19][30] , \register[19][29] , \register[19][28] ,
         \register[19][27] , \register[19][26] , \register[19][25] ,
         \register[19][24] , \register[19][23] , \register[19][22] ,
         \register[19][21] , \register[19][20] , \register[19][19] ,
         \register[19][18] , \register[19][17] , \register[19][16] ,
         \register[19][15] , \register[19][14] , \register[19][13] ,
         \register[19][12] , \register[19][11] , \register[19][10] ,
         \register[19][9] , \register[19][8] , \register[19][7] ,
         \register[19][6] , \register[19][5] , \register[19][4] ,
         \register[19][3] , \register[19][2] , \register[19][1] ,
         \register[19][0] , \register[18][31] , \register[18][30] ,
         \register[18][29] , \register[18][28] , \register[18][27] ,
         \register[18][26] , \register[18][25] , \register[18][24] ,
         \register[18][23] , \register[18][22] , \register[18][21] ,
         \register[18][20] , \register[18][19] , \register[18][18] ,
         \register[18][17] , \register[18][16] , \register[18][15] ,
         \register[18][14] , \register[18][13] , \register[18][12] ,
         \register[18][11] , \register[18][10] , \register[18][9] ,
         \register[18][8] , \register[18][7] , \register[18][6] ,
         \register[18][5] , \register[18][4] , \register[18][3] ,
         \register[18][2] , \register[18][1] , \register[18][0] ,
         \register[17][31] , \register[17][30] , \register[17][29] ,
         \register[17][28] , \register[17][27] , \register[17][26] ,
         \register[17][25] , \register[17][24] , \register[17][23] ,
         \register[17][22] , \register[17][21] , \register[17][20] ,
         \register[17][19] , \register[17][18] , \register[17][17] ,
         \register[17][16] , \register[17][15] , \register[17][14] ,
         \register[17][13] , \register[17][12] , \register[17][11] ,
         \register[17][10] , \register[17][9] , \register[17][8] ,
         \register[17][7] , \register[17][6] , \register[17][5] ,
         \register[17][4] , \register[17][3] , \register[17][2] ,
         \register[17][1] , \register[17][0] , \register[16][31] ,
         \register[16][30] , \register[16][29] , \register[16][28] ,
         \register[16][27] , \register[16][26] , \register[16][25] ,
         \register[16][24] , \register[16][23] , \register[16][22] ,
         \register[16][21] , \register[16][20] , \register[16][19] ,
         \register[16][18] , \register[16][17] , \register[16][16] ,
         \register[16][15] , \register[16][14] , \register[16][13] ,
         \register[16][12] , \register[16][11] , \register[16][10] ,
         \register[16][9] , \register[16][8] , \register[16][7] ,
         \register[16][6] , \register[16][5] , \register[16][4] ,
         \register[16][3] , \register[16][2] , \register[16][1] ,
         \register[16][0] , \register[15][31] , \register[15][30] ,
         \register[15][29] , \register[15][28] , \register[15][27] ,
         \register[15][26] , \register[15][25] , \register[15][24] ,
         \register[15][23] , \register[15][22] , \register[15][21] ,
         \register[15][20] , \register[15][19] , \register[15][18] ,
         \register[15][17] , \register[15][16] , \register[15][15] ,
         \register[15][14] , \register[15][13] , \register[15][12] ,
         \register[15][11] , \register[15][10] , \register[15][9] ,
         \register[15][8] , \register[15][7] , \register[15][6] ,
         \register[15][5] , \register[15][4] , \register[15][3] ,
         \register[15][2] , \register[15][1] , \register[15][0] ,
         \register[14][31] , \register[14][30] , \register[14][29] ,
         \register[14][28] , \register[14][27] , \register[14][26] ,
         \register[14][25] , \register[14][24] , \register[14][23] ,
         \register[14][22] , \register[14][21] , \register[14][20] ,
         \register[14][19] , \register[14][18] , \register[14][17] ,
         \register[14][16] , \register[14][15] , \register[14][14] ,
         \register[14][13] , \register[14][12] , \register[14][11] ,
         \register[14][10] , \register[14][9] , \register[14][8] ,
         \register[14][7] , \register[14][6] , \register[14][5] ,
         \register[14][4] , \register[14][3] , \register[14][2] ,
         \register[14][1] , \register[14][0] , \register[13][31] ,
         \register[13][30] , \register[13][29] , \register[13][28] ,
         \register[13][27] , \register[13][26] , \register[13][25] ,
         \register[13][24] , \register[13][23] , \register[13][22] ,
         \register[13][21] , \register[13][20] , \register[13][19] ,
         \register[13][18] , \register[13][17] , \register[13][16] ,
         \register[13][15] , \register[13][14] , \register[13][13] ,
         \register[13][12] , \register[13][11] , \register[13][10] ,
         \register[13][9] , \register[13][8] , \register[13][7] ,
         \register[13][6] , \register[13][5] , \register[13][4] ,
         \register[13][3] , \register[13][2] , \register[13][1] ,
         \register[13][0] , \register[12][31] , \register[12][30] ,
         \register[12][29] , \register[12][28] , \register[12][27] ,
         \register[12][26] , \register[12][25] , \register[12][24] ,
         \register[12][23] , \register[12][22] , \register[12][21] ,
         \register[12][20] , \register[12][19] , \register[12][18] ,
         \register[12][17] , \register[12][16] , \register[12][15] ,
         \register[12][14] , \register[12][13] , \register[12][12] ,
         \register[12][11] , \register[12][10] , \register[12][9] ,
         \register[12][8] , \register[12][7] , \register[12][6] ,
         \register[12][5] , \register[12][4] , \register[12][3] ,
         \register[12][2] , \register[12][1] , \register[12][0] ,
         \register[11][31] , \register[11][30] , \register[11][29] ,
         \register[11][28] , \register[11][27] , \register[11][26] ,
         \register[11][25] , \register[11][24] , \register[11][23] ,
         \register[11][22] , \register[11][21] , \register[11][20] ,
         \register[11][19] , \register[11][18] , \register[11][17] ,
         \register[11][16] , \register[11][15] , \register[11][14] ,
         \register[11][13] , \register[11][12] , \register[11][11] ,
         \register[11][10] , \register[11][9] , \register[11][8] ,
         \register[11][7] , \register[11][6] , \register[11][5] ,
         \register[11][4] , \register[11][3] , \register[11][2] ,
         \register[11][1] , \register[11][0] , \register[10][31] ,
         \register[10][30] , \register[10][29] , \register[10][28] ,
         \register[10][27] , \register[10][26] , \register[10][25] ,
         \register[10][24] , \register[10][23] , \register[10][22] ,
         \register[10][21] , \register[10][20] , \register[10][19] ,
         \register[10][18] , \register[10][17] , \register[10][16] ,
         \register[10][15] , \register[10][14] , \register[10][13] ,
         \register[10][12] , \register[10][11] , \register[10][10] ,
         \register[10][9] , \register[10][8] , \register[10][7] ,
         \register[10][6] , \register[10][5] , \register[10][4] ,
         \register[10][3] , \register[10][2] , \register[10][1] ,
         \register[10][0] , \register[9][31] , \register[9][30] ,
         \register[9][29] , \register[9][28] , \register[9][27] ,
         \register[9][26] , \register[9][25] , \register[9][24] ,
         \register[9][23] , \register[9][22] , \register[9][21] ,
         \register[9][20] , \register[9][19] , \register[9][18] ,
         \register[9][17] , \register[9][16] , \register[9][15] ,
         \register[9][14] , \register[9][13] , \register[9][12] ,
         \register[9][11] , \register[9][10] , \register[9][9] ,
         \register[9][8] , \register[9][7] , \register[9][6] ,
         \register[9][5] , \register[9][4] , \register[9][3] ,
         \register[9][2] , \register[9][1] , \register[9][0] ,
         \register[8][31] , \register[8][30] , \register[8][29] ,
         \register[8][28] , \register[8][27] , \register[8][26] ,
         \register[8][25] , \register[8][24] , \register[8][23] ,
         \register[8][22] , \register[8][21] , \register[8][20] ,
         \register[8][19] , \register[8][18] , \register[8][17] ,
         \register[8][16] , \register[8][15] , \register[8][14] ,
         \register[8][13] , \register[8][12] , \register[8][11] ,
         \register[8][10] , \register[8][9] , \register[8][8] ,
         \register[8][7] , \register[8][6] , \register[8][5] ,
         \register[8][4] , \register[8][3] , \register[8][2] ,
         \register[8][1] , \register[8][0] , \register[7][31] ,
         \register[7][30] , \register[7][29] , \register[7][28] ,
         \register[7][27] , \register[7][26] , \register[7][25] ,
         \register[7][24] , \register[7][23] , \register[7][22] ,
         \register[7][21] , \register[7][20] , \register[7][19] ,
         \register[7][18] , \register[7][17] , \register[7][16] ,
         \register[7][15] , \register[7][14] , \register[7][13] ,
         \register[7][12] , \register[7][11] , \register[7][10] ,
         \register[7][9] , \register[7][8] , \register[7][7] ,
         \register[7][6] , \register[7][5] , \register[7][4] ,
         \register[7][3] , \register[7][2] , \register[7][1] ,
         \register[7][0] , \register[6][31] , \register[6][30] ,
         \register[6][29] , \register[6][28] , \register[6][27] ,
         \register[6][26] , \register[6][25] , \register[6][24] ,
         \register[6][23] , \register[6][22] , \register[6][21] ,
         \register[6][20] , \register[6][19] , \register[6][18] ,
         \register[6][17] , \register[6][16] , \register[6][15] ,
         \register[6][14] , \register[6][13] , \register[6][12] ,
         \register[6][11] , \register[6][10] , \register[6][9] ,
         \register[6][8] , \register[6][7] , \register[6][6] ,
         \register[6][5] , \register[6][4] , \register[6][3] ,
         \register[6][2] , \register[6][1] , \register[6][0] ,
         \register[5][31] , \register[5][30] , \register[5][29] ,
         \register[5][28] , \register[5][27] , \register[5][26] ,
         \register[5][25] , \register[5][24] , \register[5][23] ,
         \register[5][22] , \register[5][21] , \register[5][20] ,
         \register[5][19] , \register[5][18] , \register[5][17] ,
         \register[5][16] , \register[5][15] , \register[5][14] ,
         \register[5][13] , \register[5][12] , \register[5][11] ,
         \register[5][10] , \register[5][9] , \register[5][8] ,
         \register[5][7] , \register[5][6] , \register[5][5] ,
         \register[5][4] , \register[5][3] , \register[5][2] ,
         \register[5][1] , \register[5][0] , \register[4][31] ,
         \register[4][30] , \register[4][29] , \register[4][28] ,
         \register[4][27] , \register[4][26] , \register[4][25] ,
         \register[4][24] , \register[4][23] , \register[4][22] ,
         \register[4][21] , \register[4][20] , \register[4][19] ,
         \register[4][18] , \register[4][17] , \register[4][16] ,
         \register[4][15] , \register[4][14] , \register[4][13] ,
         \register[4][12] , \register[4][11] , \register[4][10] ,
         \register[4][9] , \register[4][8] , \register[4][7] ,
         \register[4][6] , \register[4][5] , \register[4][4] ,
         \register[4][3] , \register[4][2] , \register[4][1] ,
         \register[4][0] , \register[3][31] , \register[3][30] ,
         \register[3][29] , \register[3][28] , \register[3][27] ,
         \register[3][26] , \register[3][25] , \register[3][24] ,
         \register[3][23] , \register[3][22] , \register[3][21] ,
         \register[3][20] , \register[3][19] , \register[3][18] ,
         \register[3][17] , \register[3][16] , \register[3][15] ,
         \register[3][14] , \register[3][13] , \register[3][12] ,
         \register[3][11] , \register[3][10] , \register[3][9] ,
         \register[3][8] , \register[3][7] , \register[3][6] ,
         \register[3][5] , \register[3][4] , \register[3][3] ,
         \register[3][2] , \register[3][1] , \register[3][0] ,
         \register[2][31] , \register[2][30] , \register[2][29] ,
         \register[2][28] , \register[2][27] , \register[2][26] ,
         \register[2][25] , \register[2][24] , \register[2][23] ,
         \register[2][22] , \register[2][21] , \register[2][20] ,
         \register[2][19] , \register[2][18] , \register[2][17] ,
         \register[2][16] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[1][31] ,
         \register[1][30] , \register[1][29] , \register[1][28] ,
         \register[1][27] , \register[1][26] , \register[1][25] ,
         \register[1][24] , \register[1][23] , \register[1][22] ,
         \register[1][21] , \register[1][20] , \register[1][19] ,
         \register[1][18] , \register[1][17] , \register[1][16] ,
         \register[1][15] , \register[1][14] , \register[1][13] ,
         \register[1][12] , \register[1][11] , \register[1][10] ,
         \register[1][9] , \register[1][8] , \register[1][7] ,
         \register[1][6] , \register[1][5] , \register[1][4] ,
         \register[1][3] , \register[1][2] , \register[1][1] ,
         \register[1][0] , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432;
  assign N13 = ReadReg1[0];
  assign N14 = ReadReg1[1];
  assign N15 = ReadReg1[2];
  assign N16 = ReadReg1[3];
  assign N17 = ReadReg1[4];
  assign N18 = ReadReg2[0];
  assign N19 = ReadReg2[1];
  assign N20 = ReadReg2[2];
  assign N21 = ReadReg2[3];
  assign N22 = ReadReg2[4];

  DFFRX1 \register_reg[31][31]  ( .D(n1073), .CK(clk), .RN(n2259), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n1072), .CK(clk), .RN(n2258), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n1071), .CK(clk), .RN(n2257), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n1070), .CK(clk), .RN(n2256), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n1069), .CK(clk), .RN(n2264), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n1068), .CK(clk), .RN(n2263), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n1067), .CK(clk), .RN(n2262), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n1066), .CK(clk), .RN(n2297), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n1065), .CK(clk), .RN(n2296), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n1064), .CK(clk), .RN(n2291), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n1063), .CK(clk), .RN(n2290), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n1062), .CK(clk), .RN(n2289), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n1061), .CK(clk), .RN(n2288), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n1060), .CK(clk), .RN(n2287), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n1059), .CK(clk), .RN(n2286), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n1058), .CK(clk), .RN(n2255), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n1057), .CK(clk), .RN(n2254), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n1056), .CK(clk), .RN(n2325), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n1055), .CK(clk), .RN(n2325), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n1054), .CK(clk), .RN(n2325), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n1053), .CK(clk), .RN(n2325), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n1052), .CK(clk), .RN(n2325), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n1051), .CK(clk), .RN(n2325), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n945), .CK(clk), .RN(n2317), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n944), .CK(clk), .RN(n2317), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n943), .CK(clk), .RN(n2317), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n942), .CK(clk), .RN(n2317), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n941), .CK(clk), .RN(n2317), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n940), .CK(clk), .RN(n2317), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n939), .CK(clk), .RN(n2316), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n938), .CK(clk), .RN(n2316), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n937), .CK(clk), .RN(n2316), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n936), .CK(clk), .RN(n2316), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n935), .CK(clk), .RN(n2316), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n934), .CK(clk), .RN(n2316), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n933), .CK(clk), .RN(n2316), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n932), .CK(clk), .RN(n2316), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n931), .CK(clk), .RN(n2316), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n930), .CK(clk), .RN(n2316), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n929), .CK(clk), .RN(n2316), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n928), .CK(clk), .RN(n2316), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n927), .CK(clk), .RN(n2316), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n926), .CK(clk), .RN(n2315), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n925), .CK(clk), .RN(n2315), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n924), .CK(clk), .RN(n2315), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n923), .CK(clk), .RN(n2315), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n817), .CK(clk), .RN(n2307), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n816), .CK(clk), .RN(n2307), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n815), .CK(clk), .RN(n2307), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n814), .CK(clk), .RN(n2307), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n813), .CK(clk), .RN(n2307), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n812), .CK(clk), .RN(n2307), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n811), .CK(clk), .RN(n2307), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n810), .CK(clk), .RN(n2307), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n809), .CK(clk), .RN(n2306), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n808), .CK(clk), .RN(n2306), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n807), .CK(clk), .RN(n2306), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n806), .CK(clk), .RN(n2306), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n805), .CK(clk), .RN(n2306), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n804), .CK(clk), .RN(n2306), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n803), .CK(clk), .RN(n2306), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n802), .CK(clk), .RN(n2306), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n801), .CK(clk), .RN(n2306), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n800), .CK(clk), .RN(n2306), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n799), .CK(clk), .RN(n2306), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n798), .CK(clk), .RN(n2306), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n797), .CK(clk), .RN(n2306), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n796), .CK(clk), .RN(n2305), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n795), .CK(clk), .RN(n2305), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n689), .CK(clk), .RN(n2297), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n688), .CK(clk), .RN(n2297), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n687), .CK(clk), .RN(n2297), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n686), .CK(clk), .RN(n2297), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n685), .CK(clk), .RN(n2297), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n684), .CK(clk), .RN(n2297), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n683), .CK(clk), .RN(n2297), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n682), .CK(clk), .RN(n2297), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n681), .CK(clk), .RN(n2297), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n680), .CK(clk), .RN(n2297), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n679), .CK(clk), .RN(n2296), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n678), .CK(clk), .RN(n2296), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n677), .CK(clk), .RN(n2296), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n676), .CK(clk), .RN(n2296), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n675), .CK(clk), .RN(n2296), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n674), .CK(clk), .RN(n2296), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n673), .CK(clk), .RN(n2296), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n672), .CK(clk), .RN(n2296), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n671), .CK(clk), .RN(n2296), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n670), .CK(clk), .RN(n2296), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n669), .CK(clk), .RN(n2296), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n668), .CK(clk), .RN(n2296), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n667), .CK(clk), .RN(n2296), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n561), .CK(clk), .RN(n2287), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n560), .CK(clk), .RN(n2287), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n559), .CK(clk), .RN(n2287), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n558), .CK(clk), .RN(n2287), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n557), .CK(clk), .RN(n2287), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n556), .CK(clk), .RN(n2287), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n555), .CK(clk), .RN(n2287), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n554), .CK(clk), .RN(n2287), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n553), .CK(clk), .RN(n2287), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n552), .CK(clk), .RN(n2287), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n551), .CK(clk), .RN(n2287), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n550), .CK(clk), .RN(n2287), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n549), .CK(clk), .RN(n2286), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n548), .CK(clk), .RN(n2286), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n547), .CK(clk), .RN(n2286), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n546), .CK(clk), .RN(n2286), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n545), .CK(clk), .RN(n2286), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n544), .CK(clk), .RN(n2286), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n543), .CK(clk), .RN(n2286), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n542), .CK(clk), .RN(n2286), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n541), .CK(clk), .RN(n2286), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n540), .CK(clk), .RN(n2286), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n539), .CK(clk), .RN(n2286), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n433), .CK(clk), .RN(n2278), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n432), .CK(clk), .RN(n2277), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n431), .CK(clk), .RN(n2277), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n430), .CK(clk), .RN(n2277), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n429), .CK(clk), .RN(n2277), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n428), .CK(clk), .RN(n2277), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n427), .CK(clk), .RN(n2277), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n426), .CK(clk), .RN(n2277), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n425), .CK(clk), .RN(n2277), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n424), .CK(clk), .RN(n2277), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n423), .CK(clk), .RN(n2277), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n422), .CK(clk), .RN(n2277), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n421), .CK(clk), .RN(n2277), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n420), .CK(clk), .RN(n2277), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n419), .CK(clk), .RN(n2276), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n418), .CK(clk), .RN(n2276), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n417), .CK(clk), .RN(n2276), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n416), .CK(clk), .RN(n2276), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n415), .CK(clk), .RN(n2276), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n414), .CK(clk), .RN(n2276), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n413), .CK(clk), .RN(n2276), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n412), .CK(clk), .RN(n2276), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n411), .CK(clk), .RN(n2276), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n305), .CK(clk), .RN(n2268), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n304), .CK(clk), .RN(n2268), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n303), .CK(clk), .RN(n2268), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n302), .CK(clk), .RN(n2267), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n301), .CK(clk), .RN(n2267), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n300), .CK(clk), .RN(n2267), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n299), .CK(clk), .RN(n2267), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n298), .CK(clk), .RN(n2267), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n297), .CK(clk), .RN(n2267), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n296), .CK(clk), .RN(n2267), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n295), .CK(clk), .RN(n2267), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n294), .CK(clk), .RN(n2267), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n293), .CK(clk), .RN(n2267), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n292), .CK(clk), .RN(n2267), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n291), .CK(clk), .RN(n2267), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n290), .CK(clk), .RN(n2267), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n289), .CK(clk), .RN(n2266), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n288), .CK(clk), .RN(n2266), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n287), .CK(clk), .RN(n2266), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n286), .CK(clk), .RN(n2266), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n285), .CK(clk), .RN(n2266), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n284), .CK(clk), .RN(n2266), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n283), .CK(clk), .RN(n2266), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n1009), .CK(clk), .RN(n2322), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n1008), .CK(clk), .RN(n2322), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n1007), .CK(clk), .RN(n2322), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n1006), .CK(clk), .RN(n2322), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n1005), .CK(clk), .RN(n2322), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n1004), .CK(clk), .RN(n2321), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n1003), .CK(clk), .RN(n2321), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n1002), .CK(clk), .RN(n2321), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n1001), .CK(clk), .RN(n2321), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n1000), .CK(clk), .RN(n2321), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n999), .CK(clk), .RN(n2321), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n998), .CK(clk), .RN(n2321), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n997), .CK(clk), .RN(n2321), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n996), .CK(clk), .RN(n2321), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n995), .CK(clk), .RN(n2321), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n994), .CK(clk), .RN(n2321), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n993), .CK(clk), .RN(n2321), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n992), .CK(clk), .RN(n2321), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n991), .CK(clk), .RN(n2320), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n990), .CK(clk), .RN(n2320), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n989), .CK(clk), .RN(n2320), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n988), .CK(clk), .RN(n2320), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n987), .CK(clk), .RN(n2320), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n881), .CK(clk), .RN(n2312), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n880), .CK(clk), .RN(n2312), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n879), .CK(clk), .RN(n2312), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n878), .CK(clk), .RN(n2312), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n877), .CK(clk), .RN(n2312), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n876), .CK(clk), .RN(n2312), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n875), .CK(clk), .RN(n2312), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n874), .CK(clk), .RN(n2311), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n873), .CK(clk), .RN(n2311), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n872), .CK(clk), .RN(n2311), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n871), .CK(clk), .RN(n2311), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n870), .CK(clk), .RN(n2311), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n869), .CK(clk), .RN(n2311), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n868), .CK(clk), .RN(n2311), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n867), .CK(clk), .RN(n2311), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n866), .CK(clk), .RN(n2311), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n865), .CK(clk), .RN(n2311), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n864), .CK(clk), .RN(n2311), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n863), .CK(clk), .RN(n2311), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n862), .CK(clk), .RN(n2311), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n861), .CK(clk), .RN(n2310), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n860), .CK(clk), .RN(n2310), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n859), .CK(clk), .RN(n2310), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n753), .CK(clk), .RN(n2302), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n752), .CK(clk), .RN(n2302), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n751), .CK(clk), .RN(n2302), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n750), .CK(clk), .RN(n2302), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n749), .CK(clk), .RN(n2302), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n748), .CK(clk), .RN(n2302), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n747), .CK(clk), .RN(n2302), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n746), .CK(clk), .RN(n2302), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n745), .CK(clk), .RN(n2302), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n744), .CK(clk), .RN(n2301), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n743), .CK(clk), .RN(n2301), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n742), .CK(clk), .RN(n2301), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n741), .CK(clk), .RN(n2301), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n740), .CK(clk), .RN(n2301), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n739), .CK(clk), .RN(n2301), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n738), .CK(clk), .RN(n2301), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n737), .CK(clk), .RN(n2301), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n736), .CK(clk), .RN(n2301), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n735), .CK(clk), .RN(n2301), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n734), .CK(clk), .RN(n2301), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n733), .CK(clk), .RN(n2301), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n732), .CK(clk), .RN(n2301), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n731), .CK(clk), .RN(n2300), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n625), .CK(clk), .RN(n2292), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n624), .CK(clk), .RN(n2292), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n623), .CK(clk), .RN(n2292), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n622), .CK(clk), .RN(n2292), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n621), .CK(clk), .RN(n2292), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n620), .CK(clk), .RN(n2292), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n619), .CK(clk), .RN(n2292), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n618), .CK(clk), .RN(n2292), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n617), .CK(clk), .RN(n2292), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n616), .CK(clk), .RN(n2292), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n615), .CK(clk), .RN(n2292), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n614), .CK(clk), .RN(n2291), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n613), .CK(clk), .RN(n2291), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n612), .CK(clk), .RN(n2291), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n611), .CK(clk), .RN(n2291), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n610), .CK(clk), .RN(n2291), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n609), .CK(clk), .RN(n2291), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n608), .CK(clk), .RN(n2291), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n607), .CK(clk), .RN(n2291), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n606), .CK(clk), .RN(n2291), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n605), .CK(clk), .RN(n2291), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n604), .CK(clk), .RN(n2291), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n603), .CK(clk), .RN(n2291), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n497), .CK(clk), .RN(n2282), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n496), .CK(clk), .RN(n2282), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n495), .CK(clk), .RN(n2282), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n494), .CK(clk), .RN(n2282), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n493), .CK(clk), .RN(n2282), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n492), .CK(clk), .RN(n2282), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n491), .CK(clk), .RN(n2282), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n490), .CK(clk), .RN(n2282), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n489), .CK(clk), .RN(n2282), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n488), .CK(clk), .RN(n2282), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n487), .CK(clk), .RN(n2282), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n486), .CK(clk), .RN(n2282), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n485), .CK(clk), .RN(n2282), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n484), .CK(clk), .RN(n2281), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n483), .CK(clk), .RN(n2281), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n482), .CK(clk), .RN(n2281), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n481), .CK(clk), .RN(n2281), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n480), .CK(clk), .RN(n2281), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n479), .CK(clk), .RN(n2281), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n478), .CK(clk), .RN(n2281), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n477), .CK(clk), .RN(n2281), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n476), .CK(clk), .RN(n2281), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n475), .CK(clk), .RN(n2281), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n369), .CK(clk), .RN(n2273), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n368), .CK(clk), .RN(n2273), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n367), .CK(clk), .RN(n2272), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n366), .CK(clk), .RN(n2272), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n365), .CK(clk), .RN(n2272), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n364), .CK(clk), .RN(n2272), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n363), .CK(clk), .RN(n2272), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n362), .CK(clk), .RN(n2272), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n361), .CK(clk), .RN(n2272), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n360), .CK(clk), .RN(n2272), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n359), .CK(clk), .RN(n2272), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n358), .CK(clk), .RN(n2272), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n357), .CK(clk), .RN(n2272), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n356), .CK(clk), .RN(n2272), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n355), .CK(clk), .RN(n2272), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n354), .CK(clk), .RN(n2271), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n353), .CK(clk), .RN(n2271), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n352), .CK(clk), .RN(n2271), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n351), .CK(clk), .RN(n2271), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n350), .CK(clk), .RN(n2271), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n349), .CK(clk), .RN(n2271), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n348), .CK(clk), .RN(n2271), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n347), .CK(clk), .RN(n2271), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n241), .CK(clk), .RN(n2263), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n240), .CK(clk), .RN(n2263), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n239), .CK(clk), .RN(n2263), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n238), .CK(clk), .RN(n2263), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n237), .CK(clk), .RN(n2262), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n236), .CK(clk), .RN(n2262), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n235), .CK(clk), .RN(n2262), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n234), .CK(clk), .RN(n2262), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n233), .CK(clk), .RN(n2262), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n232), .CK(clk), .RN(n2262), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n231), .CK(clk), .RN(n2262), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n230), .CK(clk), .RN(n2262), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n229), .CK(clk), .RN(n2262), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n228), .CK(clk), .RN(n2262), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n227), .CK(clk), .RN(n2262), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n226), .CK(clk), .RN(n2262), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n225), .CK(clk), .RN(n2262), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n224), .CK(clk), .RN(n2261), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n223), .CK(clk), .RN(n2261), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n222), .CK(clk), .RN(n2261), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n221), .CK(clk), .RN(n2261), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n220), .CK(clk), .RN(n2261), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n219), .CK(clk), .RN(n2261), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n977), .CK(clk), .RN(n2319), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n976), .CK(clk), .RN(n2319), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n975), .CK(clk), .RN(n2319), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n974), .CK(clk), .RN(n2319), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n973), .CK(clk), .RN(n2319), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n972), .CK(clk), .RN(n2319), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n971), .CK(clk), .RN(n2319), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n970), .CK(clk), .RN(n2319), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n969), .CK(clk), .RN(n2319), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n968), .CK(clk), .RN(n2319), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n967), .CK(clk), .RN(n2319), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n966), .CK(clk), .RN(n2319), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n965), .CK(clk), .RN(n2318), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n964), .CK(clk), .RN(n2318), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n963), .CK(clk), .RN(n2318), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n962), .CK(clk), .RN(n2318), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n961), .CK(clk), .RN(n2318), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n960), .CK(clk), .RN(n2318), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n959), .CK(clk), .RN(n2318), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n958), .CK(clk), .RN(n2318), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n957), .CK(clk), .RN(n2318), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n956), .CK(clk), .RN(n2318), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n955), .CK(clk), .RN(n2318), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n849), .CK(clk), .RN(n2310), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n848), .CK(clk), .RN(n2309), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n847), .CK(clk), .RN(n2309), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n846), .CK(clk), .RN(n2309), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n845), .CK(clk), .RN(n2309), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n844), .CK(clk), .RN(n2309), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n843), .CK(clk), .RN(n2309), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n842), .CK(clk), .RN(n2309), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n841), .CK(clk), .RN(n2309), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n840), .CK(clk), .RN(n2309), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n839), .CK(clk), .RN(n2309), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n838), .CK(clk), .RN(n2309), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n837), .CK(clk), .RN(n2309), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n836), .CK(clk), .RN(n2309), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n835), .CK(clk), .RN(n2308), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n834), .CK(clk), .RN(n2308), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n833), .CK(clk), .RN(n2308), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n832), .CK(clk), .RN(n2308), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n831), .CK(clk), .RN(n2308), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n830), .CK(clk), .RN(n2308), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n829), .CK(clk), .RN(n2308), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n828), .CK(clk), .RN(n2308), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n827), .CK(clk), .RN(n2308), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n721), .CK(clk), .RN(n2300), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n720), .CK(clk), .RN(n2300), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n719), .CK(clk), .RN(n2300), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n718), .CK(clk), .RN(n2299), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n717), .CK(clk), .RN(n2299), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n716), .CK(clk), .RN(n2299), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n715), .CK(clk), .RN(n2299), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n714), .CK(clk), .RN(n2299), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n713), .CK(clk), .RN(n2299), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n712), .CK(clk), .RN(n2299), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n711), .CK(clk), .RN(n2299), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n710), .CK(clk), .RN(n2299), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n709), .CK(clk), .RN(n2299), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n708), .CK(clk), .RN(n2299), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n707), .CK(clk), .RN(n2299), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n706), .CK(clk), .RN(n2299), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n705), .CK(clk), .RN(n2298), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n704), .CK(clk), .RN(n2298), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n703), .CK(clk), .RN(n2298), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n702), .CK(clk), .RN(n2298), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n701), .CK(clk), .RN(n2298), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n700), .CK(clk), .RN(n2298), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n699), .CK(clk), .RN(n2298), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n593), .CK(clk), .RN(n2290), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n592), .CK(clk), .RN(n2290), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n591), .CK(clk), .RN(n2290), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n590), .CK(clk), .RN(n2290), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n589), .CK(clk), .RN(n2290), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n588), .CK(clk), .RN(n2289), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n587), .CK(clk), .RN(n2289), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n586), .CK(clk), .RN(n2289), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n585), .CK(clk), .RN(n2289), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n584), .CK(clk), .RN(n2289), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n583), .CK(clk), .RN(n2289), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n582), .CK(clk), .RN(n2289), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n581), .CK(clk), .RN(n2289), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n580), .CK(clk), .RN(n2289), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n579), .CK(clk), .RN(n2289), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n578), .CK(clk), .RN(n2289), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n577), .CK(clk), .RN(n2289), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n576), .CK(clk), .RN(n2289), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n575), .CK(clk), .RN(n2288), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n574), .CK(clk), .RN(n2288), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n573), .CK(clk), .RN(n2288), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n572), .CK(clk), .RN(n2288), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n571), .CK(clk), .RN(n2288), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n465), .CK(clk), .RN(n2280), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n464), .CK(clk), .RN(n2280), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n463), .CK(clk), .RN(n2280), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n462), .CK(clk), .RN(n2280), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n461), .CK(clk), .RN(n2280), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n460), .CK(clk), .RN(n2280), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n459), .CK(clk), .RN(n2280), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n458), .CK(clk), .RN(n2279), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n457), .CK(clk), .RN(n2279), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n456), .CK(clk), .RN(n2279), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n455), .CK(clk), .RN(n2279), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n454), .CK(clk), .RN(n2279), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n453), .CK(clk), .RN(n2279), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n452), .CK(clk), .RN(n2279), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n451), .CK(clk), .RN(n2279), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n450), .CK(clk), .RN(n2279), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n449), .CK(clk), .RN(n2279), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n448), .CK(clk), .RN(n2279), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n447), .CK(clk), .RN(n2279), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n446), .CK(clk), .RN(n2279), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n445), .CK(clk), .RN(n2278), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n444), .CK(clk), .RN(n2278), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n443), .CK(clk), .RN(n2278), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n337), .CK(clk), .RN(n2270), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n336), .CK(clk), .RN(n2270), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n335), .CK(clk), .RN(n2270), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n334), .CK(clk), .RN(n2270), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n333), .CK(clk), .RN(n2270), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n332), .CK(clk), .RN(n2270), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n331), .CK(clk), .RN(n2270), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n330), .CK(clk), .RN(n2270), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n329), .CK(clk), .RN(n2270), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n328), .CK(clk), .RN(n2269), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n327), .CK(clk), .RN(n2269), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n326), .CK(clk), .RN(n2269), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n325), .CK(clk), .RN(n2269), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n324), .CK(clk), .RN(n2269), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n323), .CK(clk), .RN(n2269), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n322), .CK(clk), .RN(n2269), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n321), .CK(clk), .RN(n2269), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n320), .CK(clk), .RN(n2269), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n319), .CK(clk), .RN(n2269), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n318), .CK(clk), .RN(n2269), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n317), .CK(clk), .RN(n2269), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n316), .CK(clk), .RN(n2269), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n315), .CK(clk), .RN(n2268), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n209), .CK(clk), .RN(n2260), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n208), .CK(clk), .RN(n2260), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n207), .CK(clk), .RN(n2260), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n206), .CK(clk), .RN(n2260), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n205), .CK(clk), .RN(n2260), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n204), .CK(clk), .RN(n2260), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n203), .CK(clk), .RN(n2260), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n202), .CK(clk), .RN(n2260), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n201), .CK(clk), .RN(n2260), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n200), .CK(clk), .RN(n2260), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n199), .CK(clk), .RN(n2260), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n198), .CK(clk), .RN(n2259), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n197), .CK(clk), .RN(n2259), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n196), .CK(clk), .RN(n2259), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n195), .CK(clk), .RN(n2259), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n194), .CK(clk), .RN(n2259), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n193), .CK(clk), .RN(n2259), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n192), .CK(clk), .RN(n2259), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n191), .CK(clk), .RN(n2259), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n190), .CK(clk), .RN(n2259), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n189), .CK(clk), .RN(n2259), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n188), .CK(clk), .RN(n2259), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n187), .CK(clk), .RN(n2259), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n1041), .CK(clk), .RN(n2324), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n1040), .CK(clk), .RN(n2324), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n1039), .CK(clk), .RN(n2324), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n1038), .CK(clk), .RN(n2324), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n1037), .CK(clk), .RN(n2324), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n1036), .CK(clk), .RN(n2324), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n1035), .CK(clk), .RN(n2324), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n1034), .CK(clk), .RN(n2324), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n1033), .CK(clk), .RN(n2324), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n1032), .CK(clk), .RN(n2324), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n1031), .CK(clk), .RN(n2324), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n1030), .CK(clk), .RN(n2323), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n1029), .CK(clk), .RN(n2323), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n1028), .CK(clk), .RN(n2323), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n1027), .CK(clk), .RN(n2323), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n1026), .CK(clk), .RN(n2323), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n1025), .CK(clk), .RN(n2323), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n1024), .CK(clk), .RN(n2323), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n1023), .CK(clk), .RN(n2323), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n1022), .CK(clk), .RN(n2323), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n1021), .CK(clk), .RN(n2323), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n1020), .CK(clk), .RN(n2323), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n1019), .CK(clk), .RN(n2323), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n913), .CK(clk), .RN(n2314), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n912), .CK(clk), .RN(n2314), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n911), .CK(clk), .RN(n2314), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n910), .CK(clk), .RN(n2314), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n909), .CK(clk), .RN(n2314), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n908), .CK(clk), .RN(n2314), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n907), .CK(clk), .RN(n2314), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n906), .CK(clk), .RN(n2314), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n905), .CK(clk), .RN(n2314), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n904), .CK(clk), .RN(n2314), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n903), .CK(clk), .RN(n2314), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n902), .CK(clk), .RN(n2314), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n901), .CK(clk), .RN(n2314), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n900), .CK(clk), .RN(n2313), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n899), .CK(clk), .RN(n2313), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n898), .CK(clk), .RN(n2313), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n897), .CK(clk), .RN(n2313), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n896), .CK(clk), .RN(n2313), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n895), .CK(clk), .RN(n2313), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n894), .CK(clk), .RN(n2313), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n893), .CK(clk), .RN(n2313), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n892), .CK(clk), .RN(n2313), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n891), .CK(clk), .RN(n2313), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n785), .CK(clk), .RN(n2305), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n784), .CK(clk), .RN(n2305), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n783), .CK(clk), .RN(n2304), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n782), .CK(clk), .RN(n2304), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n781), .CK(clk), .RN(n2304), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n780), .CK(clk), .RN(n2304), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n779), .CK(clk), .RN(n2304), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n778), .CK(clk), .RN(n2304), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n777), .CK(clk), .RN(n2304), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n776), .CK(clk), .RN(n2304), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n775), .CK(clk), .RN(n2304), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n774), .CK(clk), .RN(n2304), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n773), .CK(clk), .RN(n2304), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n772), .CK(clk), .RN(n2304), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n771), .CK(clk), .RN(n2304), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n770), .CK(clk), .RN(n2303), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n769), .CK(clk), .RN(n2303), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n768), .CK(clk), .RN(n2303), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n767), .CK(clk), .RN(n2303), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n766), .CK(clk), .RN(n2303), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n765), .CK(clk), .RN(n2303), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n764), .CK(clk), .RN(n2303), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n763), .CK(clk), .RN(n2303), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n657), .CK(clk), .RN(n2295), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n656), .CK(clk), .RN(n2295), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n655), .CK(clk), .RN(n2295), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n654), .CK(clk), .RN(n2295), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n653), .CK(clk), .RN(n2294), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n652), .CK(clk), .RN(n2294), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n651), .CK(clk), .RN(n2294), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n650), .CK(clk), .RN(n2294), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n649), .CK(clk), .RN(n2294), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n648), .CK(clk), .RN(n2294), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n647), .CK(clk), .RN(n2294), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n646), .CK(clk), .RN(n2294), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n645), .CK(clk), .RN(n2294), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n644), .CK(clk), .RN(n2294), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n643), .CK(clk), .RN(n2294), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n642), .CK(clk), .RN(n2294), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n641), .CK(clk), .RN(n2294), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n640), .CK(clk), .RN(n2293), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n639), .CK(clk), .RN(n2293), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n638), .CK(clk), .RN(n2293), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n637), .CK(clk), .RN(n2293), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n636), .CK(clk), .RN(n2293), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n635), .CK(clk), .RN(n2293), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n529), .CK(clk), .RN(n2285), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n528), .CK(clk), .RN(n2285), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n527), .CK(clk), .RN(n2285), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n526), .CK(clk), .RN(n2285), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n525), .CK(clk), .RN(n2285), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n524), .CK(clk), .RN(n2285), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n523), .CK(clk), .RN(n2284), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n522), .CK(clk), .RN(n2284), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n521), .CK(clk), .RN(n2284), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n520), .CK(clk), .RN(n2284), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n519), .CK(clk), .RN(n2284), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n518), .CK(clk), .RN(n2284), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n517), .CK(clk), .RN(n2284), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n516), .CK(clk), .RN(n2284), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n515), .CK(clk), .RN(n2284), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n514), .CK(clk), .RN(n2284), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n513), .CK(clk), .RN(n2284), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n512), .CK(clk), .RN(n2284), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n511), .CK(clk), .RN(n2284), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n510), .CK(clk), .RN(n2283), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n509), .CK(clk), .RN(n2283), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n508), .CK(clk), .RN(n2283), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n507), .CK(clk), .RN(n2283), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n401), .CK(clk), .RN(n2275), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n400), .CK(clk), .RN(n2275), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n399), .CK(clk), .RN(n2275), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n398), .CK(clk), .RN(n2275), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n397), .CK(clk), .RN(n2275), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n396), .CK(clk), .RN(n2275), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n395), .CK(clk), .RN(n2275), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n394), .CK(clk), .RN(n2275), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n393), .CK(clk), .RN(n2274), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n392), .CK(clk), .RN(n2274), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n391), .CK(clk), .RN(n2274), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n390), .CK(clk), .RN(n2274), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n389), .CK(clk), .RN(n2274), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n388), .CK(clk), .RN(n2274), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n387), .CK(clk), .RN(n2274), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n386), .CK(clk), .RN(n2274), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n385), .CK(clk), .RN(n2274), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n384), .CK(clk), .RN(n2274), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n383), .CK(clk), .RN(n2274), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n382), .CK(clk), .RN(n2274), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n381), .CK(clk), .RN(n2274), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n380), .CK(clk), .RN(n2273), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n379), .CK(clk), .RN(n2273), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n273), .CK(clk), .RN(n2265), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n272), .CK(clk), .RN(n2265), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n271), .CK(clk), .RN(n2265), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n270), .CK(clk), .RN(n2265), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n269), .CK(clk), .RN(n2265), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n268), .CK(clk), .RN(n2265), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n267), .CK(clk), .RN(n2265), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n266), .CK(clk), .RN(n2265), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n265), .CK(clk), .RN(n2265), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n264), .CK(clk), .RN(n2265), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n263), .CK(clk), .RN(n2264), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n262), .CK(clk), .RN(n2264), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n261), .CK(clk), .RN(n2264), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n260), .CK(clk), .RN(n2264), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n259), .CK(clk), .RN(n2264), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n258), .CK(clk), .RN(n2264), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n257), .CK(clk), .RN(n2264), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n256), .CK(clk), .RN(n2264), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n255), .CK(clk), .RN(n2264), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n254), .CK(clk), .RN(n2264), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n253), .CK(clk), .RN(n2264), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n252), .CK(clk), .RN(n2264), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n251), .CK(clk), .RN(n2264), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[3][31]  ( .D(n177), .CK(clk), .RN(n2258), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n176), .CK(clk), .RN(n2258), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n175), .CK(clk), .RN(n2258), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n174), .CK(clk), .RN(n2258), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n173), .CK(clk), .RN(n2258), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n172), .CK(clk), .RN(n2257), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n171), .CK(clk), .RN(n2257), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n170), .CK(clk), .RN(n2257), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n169), .CK(clk), .RN(n2257), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n168), .CK(clk), .RN(n2257), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n167), .CK(clk), .RN(n2257), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n166), .CK(clk), .RN(n2257), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n165), .CK(clk), .RN(n2257), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n164), .CK(clk), .RN(n2257), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n163), .CK(clk), .RN(n2257), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n162), .CK(clk), .RN(n2257), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n161), .CK(clk), .RN(n2257), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n160), .CK(clk), .RN(n2257), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n159), .CK(clk), .RN(n2256), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n158), .CK(clk), .RN(n2256), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n157), .CK(clk), .RN(n2256), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n156), .CK(clk), .RN(n2256), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n155), .CK(clk), .RN(n2256), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n113), .CK(clk), .RN(n2295), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n112), .CK(clk), .RN(n2294), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n111), .CK(clk), .RN(n2293), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n110), .CK(clk), .RN(n2292), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n109), .CK(clk), .RN(n2261), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n108), .CK(clk), .RN(n2260), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n107), .CK(clk), .RN(n2255), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n106), .CK(clk), .RN(n2255), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n105), .CK(clk), .RN(n2255), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n104), .CK(clk), .RN(n2255), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n103), .CK(clk), .RN(n2255), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n102), .CK(clk), .RN(n2255), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n101), .CK(clk), .RN(n2255), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n100), .CK(clk), .RN(n2255), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n99), .CK(clk), .RN(n2255), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n98), .CK(clk), .RN(n2255), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n97), .CK(clk), .RN(n2255), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n96), .CK(clk), .RN(n2255), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n95), .CK(clk), .RN(n2255), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n94), .CK(clk), .RN(n2254), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n93), .CK(clk), .RN(n2254), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n92), .CK(clk), .RN(n2254), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n91), .CK(clk), .RN(n2254), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n1050), .CK(clk), .RN(n2325), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n1049), .CK(clk), .RN(n2325), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n1048), .CK(clk), .RN(n2325), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n1047), .CK(clk), .RN(n2325), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n1046), .CK(clk), .RN(n2325), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n1045), .CK(clk), .RN(n2325), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n1044), .CK(clk), .RN(n2325), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n1043), .CK(clk), .RN(n2324), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n1042), .CK(clk), .RN(n2324), .Q(
        \register[31][0] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n922), .CK(clk), .RN(n2315), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n921), .CK(clk), .RN(n2315), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n920), .CK(clk), .RN(n2315), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n919), .CK(clk), .RN(n2315), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n918), .CK(clk), .RN(n2315), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n917), .CK(clk), .RN(n2315), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n916), .CK(clk), .RN(n2315), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n915), .CK(clk), .RN(n2315), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n914), .CK(clk), .RN(n2315), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n794), .CK(clk), .RN(n2305), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n793), .CK(clk), .RN(n2305), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n792), .CK(clk), .RN(n2305), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n791), .CK(clk), .RN(n2305), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n790), .CK(clk), .RN(n2305), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n789), .CK(clk), .RN(n2305), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n788), .CK(clk), .RN(n2305), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n787), .CK(clk), .RN(n2305), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n786), .CK(clk), .RN(n2305), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n666), .CK(clk), .RN(n2295), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n665), .CK(clk), .RN(n2295), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n664), .CK(clk), .RN(n2295), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n663), .CK(clk), .RN(n2295), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n662), .CK(clk), .RN(n2295), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n661), .CK(clk), .RN(n2295), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n660), .CK(clk), .RN(n2295), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n659), .CK(clk), .RN(n2295), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n658), .CK(clk), .RN(n2295), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n538), .CK(clk), .RN(n2286), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n537), .CK(clk), .RN(n2286), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n536), .CK(clk), .RN(n2285), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n535), .CK(clk), .RN(n2285), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n534), .CK(clk), .RN(n2285), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n533), .CK(clk), .RN(n2285), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n532), .CK(clk), .RN(n2285), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n531), .CK(clk), .RN(n2285), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n530), .CK(clk), .RN(n2285), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n410), .CK(clk), .RN(n2276), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n409), .CK(clk), .RN(n2276), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n408), .CK(clk), .RN(n2276), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n407), .CK(clk), .RN(n2276), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n406), .CK(clk), .RN(n2275), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n405), .CK(clk), .RN(n2275), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n404), .CK(clk), .RN(n2275), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n403), .CK(clk), .RN(n2275), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n402), .CK(clk), .RN(n2275), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n282), .CK(clk), .RN(n2266), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n281), .CK(clk), .RN(n2266), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n280), .CK(clk), .RN(n2266), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n279), .CK(clk), .RN(n2266), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n278), .CK(clk), .RN(n2266), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n277), .CK(clk), .RN(n2266), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n276), .CK(clk), .RN(n2265), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n275), .CK(clk), .RN(n2265), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n274), .CK(clk), .RN(n2265), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n986), .CK(clk), .RN(n2320), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n985), .CK(clk), .RN(n2320), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n984), .CK(clk), .RN(n2320), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n983), .CK(clk), .RN(n2320), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n982), .CK(clk), .RN(n2320), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n981), .CK(clk), .RN(n2320), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n980), .CK(clk), .RN(n2320), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n979), .CK(clk), .RN(n2320), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n978), .CK(clk), .RN(n2319), .Q(
        \register[29][0] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n858), .CK(clk), .RN(n2310), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n857), .CK(clk), .RN(n2310), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n856), .CK(clk), .RN(n2310), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n855), .CK(clk), .RN(n2310), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n854), .CK(clk), .RN(n2310), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n853), .CK(clk), .RN(n2310), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n852), .CK(clk), .RN(n2310), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n851), .CK(clk), .RN(n2310), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n850), .CK(clk), .RN(n2310), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n730), .CK(clk), .RN(n2300), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n729), .CK(clk), .RN(n2300), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n728), .CK(clk), .RN(n2300), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n727), .CK(clk), .RN(n2300), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n726), .CK(clk), .RN(n2300), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n725), .CK(clk), .RN(n2300), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n724), .CK(clk), .RN(n2300), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n723), .CK(clk), .RN(n2300), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n722), .CK(clk), .RN(n2300), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n602), .CK(clk), .RN(n2291), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n601), .CK(clk), .RN(n2290), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n600), .CK(clk), .RN(n2290), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n599), .CK(clk), .RN(n2290), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n598), .CK(clk), .RN(n2290), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n597), .CK(clk), .RN(n2290), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n596), .CK(clk), .RN(n2290), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n595), .CK(clk), .RN(n2290), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n594), .CK(clk), .RN(n2290), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n474), .CK(clk), .RN(n2281), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n473), .CK(clk), .RN(n2281), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n472), .CK(clk), .RN(n2281), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n471), .CK(clk), .RN(n2280), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n470), .CK(clk), .RN(n2280), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n469), .CK(clk), .RN(n2280), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n468), .CK(clk), .RN(n2280), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n467), .CK(clk), .RN(n2280), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n466), .CK(clk), .RN(n2280), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n346), .CK(clk), .RN(n2271), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n345), .CK(clk), .RN(n2271), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n344), .CK(clk), .RN(n2271), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n343), .CK(clk), .RN(n2271), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n342), .CK(clk), .RN(n2271), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n341), .CK(clk), .RN(n2270), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n340), .CK(clk), .RN(n2270), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n339), .CK(clk), .RN(n2270), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n338), .CK(clk), .RN(n2270), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n218), .CK(clk), .RN(n2261), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n217), .CK(clk), .RN(n2261), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n216), .CK(clk), .RN(n2261), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n215), .CK(clk), .RN(n2261), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n214), .CK(clk), .RN(n2261), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n213), .CK(clk), .RN(n2261), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n212), .CK(clk), .RN(n2261), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n211), .CK(clk), .RN(n2260), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n210), .CK(clk), .RN(n2260), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n954), .CK(clk), .RN(n2318), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n953), .CK(clk), .RN(n2318), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n952), .CK(clk), .RN(n2317), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n951), .CK(clk), .RN(n2317), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n950), .CK(clk), .RN(n2317), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n949), .CK(clk), .RN(n2317), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n948), .CK(clk), .RN(n2317), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n947), .CK(clk), .RN(n2317), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][0]  ( .D(n946), .CK(clk), .RN(n2317), .Q(
        \register[28][0] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n826), .CK(clk), .RN(n2308), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n825), .CK(clk), .RN(n2308), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n824), .CK(clk), .RN(n2308), .Q(
        \register[24][6] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n823), .CK(clk), .RN(n2308), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n822), .CK(clk), .RN(n2307), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n821), .CK(clk), .RN(n2307), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n820), .CK(clk), .RN(n2307), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n819), .CK(clk), .RN(n2307), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n818), .CK(clk), .RN(n2307), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n698), .CK(clk), .RN(n2298), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n697), .CK(clk), .RN(n2298), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n696), .CK(clk), .RN(n2298), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n695), .CK(clk), .RN(n2298), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n694), .CK(clk), .RN(n2298), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n693), .CK(clk), .RN(n2298), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n692), .CK(clk), .RN(n2297), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n691), .CK(clk), .RN(n2297), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[20][0]  ( .D(n690), .CK(clk), .RN(n2297), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n570), .CK(clk), .RN(n2288), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n569), .CK(clk), .RN(n2288), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n568), .CK(clk), .RN(n2288), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n567), .CK(clk), .RN(n2288), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n566), .CK(clk), .RN(n2288), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n565), .CK(clk), .RN(n2288), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n564), .CK(clk), .RN(n2288), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n563), .CK(clk), .RN(n2288), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n562), .CK(clk), .RN(n2287), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n442), .CK(clk), .RN(n2278), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n441), .CK(clk), .RN(n2278), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n440), .CK(clk), .RN(n2278), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n439), .CK(clk), .RN(n2278), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n438), .CK(clk), .RN(n2278), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n437), .CK(clk), .RN(n2278), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n436), .CK(clk), .RN(n2278), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n435), .CK(clk), .RN(n2278), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n434), .CK(clk), .RN(n2278), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n314), .CK(clk), .RN(n2268), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n313), .CK(clk), .RN(n2268), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n312), .CK(clk), .RN(n2268), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n311), .CK(clk), .RN(n2268), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n310), .CK(clk), .RN(n2268), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n309), .CK(clk), .RN(n2268), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n308), .CK(clk), .RN(n2268), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n307), .CK(clk), .RN(n2268), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n306), .CK(clk), .RN(n2268), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n186), .CK(clk), .RN(n2259), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n185), .CK(clk), .RN(n2258), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n184), .CK(clk), .RN(n2258), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n183), .CK(clk), .RN(n2258), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n182), .CK(clk), .RN(n2258), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n181), .CK(clk), .RN(n2258), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n180), .CK(clk), .RN(n2258), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n179), .CK(clk), .RN(n2258), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n178), .CK(clk), .RN(n2258), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n1018), .CK(clk), .RN(n2323), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n1017), .CK(clk), .RN(n2322), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n1016), .CK(clk), .RN(n2322), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n1015), .CK(clk), .RN(n2322), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n1014), .CK(clk), .RN(n2322), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n1013), .CK(clk), .RN(n2322), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n1012), .CK(clk), .RN(n2322), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n1011), .CK(clk), .RN(n2322), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][0]  ( .D(n1010), .CK(clk), .RN(n2322), .Q(
        \register[30][0] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n890), .CK(clk), .RN(n2313), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n889), .CK(clk), .RN(n2313), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n888), .CK(clk), .RN(n2313), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n887), .CK(clk), .RN(n2312), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n886), .CK(clk), .RN(n2312), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n885), .CK(clk), .RN(n2312), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n884), .CK(clk), .RN(n2312), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n883), .CK(clk), .RN(n2312), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n882), .CK(clk), .RN(n2312), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n762), .CK(clk), .RN(n2303), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n761), .CK(clk), .RN(n2303), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n760), .CK(clk), .RN(n2303), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n759), .CK(clk), .RN(n2303), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n758), .CK(clk), .RN(n2303), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n757), .CK(clk), .RN(n2302), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n756), .CK(clk), .RN(n2302), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n755), .CK(clk), .RN(n2302), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n754), .CK(clk), .RN(n2302), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n634), .CK(clk), .RN(n2293), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n633), .CK(clk), .RN(n2293), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n632), .CK(clk), .RN(n2293), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n631), .CK(clk), .RN(n2293), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n630), .CK(clk), .RN(n2293), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n629), .CK(clk), .RN(n2293), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n628), .CK(clk), .RN(n2293), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n627), .CK(clk), .RN(n2292), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n626), .CK(clk), .RN(n2292), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n506), .CK(clk), .RN(n2283), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n505), .CK(clk), .RN(n2283), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n504), .CK(clk), .RN(n2283), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n503), .CK(clk), .RN(n2283), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n502), .CK(clk), .RN(n2283), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n501), .CK(clk), .RN(n2283), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n500), .CK(clk), .RN(n2283), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n499), .CK(clk), .RN(n2283), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n498), .CK(clk), .RN(n2283), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n378), .CK(clk), .RN(n2273), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n377), .CK(clk), .RN(n2273), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n376), .CK(clk), .RN(n2273), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n375), .CK(clk), .RN(n2273), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n374), .CK(clk), .RN(n2273), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n373), .CK(clk), .RN(n2273), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n372), .CK(clk), .RN(n2273), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n371), .CK(clk), .RN(n2273), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n370), .CK(clk), .RN(n2273), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n250), .CK(clk), .RN(n2263), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n249), .CK(clk), .RN(n2263), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n248), .CK(clk), .RN(n2263), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n247), .CK(clk), .RN(n2263), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n246), .CK(clk), .RN(n2263), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n245), .CK(clk), .RN(n2263), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n244), .CK(clk), .RN(n2263), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n243), .CK(clk), .RN(n2263), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n242), .CK(clk), .RN(n2263), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n154), .CK(clk), .RN(n2256), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n153), .CK(clk), .RN(n2256), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n152), .CK(clk), .RN(n2256), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n151), .CK(clk), .RN(n2256), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n150), .CK(clk), .RN(n2256), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n149), .CK(clk), .RN(n2256), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n148), .CK(clk), .RN(n2256), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n147), .CK(clk), .RN(n2256), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n146), .CK(clk), .RN(n2254), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n90), .CK(clk), .RN(n2254), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n89), .CK(clk), .RN(n2254), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n88), .CK(clk), .RN(n2254), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n87), .CK(clk), .RN(n2254), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n86), .CK(clk), .RN(n2254), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n85), .CK(clk), .RN(n2254), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n84), .CK(clk), .RN(n2254), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n82), .CK(clk), .RN(n2254), .Q(
        \register[1][0] ) );
  DFFRX1 \register_reg[2][31]  ( .D(n145), .CK(clk), .RN(n2253), .Q(
        \register[2][31] ), .QN(n2396) );
  DFFRX1 \register_reg[2][30]  ( .D(n144), .CK(clk), .RN(n2253), .Q(
        \register[2][30] ), .QN(n2395) );
  DFFRX1 \register_reg[2][29]  ( .D(n143), .CK(clk), .RN(n2253), .Q(
        \register[2][29] ), .QN(n2394) );
  DFFRX1 \register_reg[2][28]  ( .D(n142), .CK(clk), .RN(n2253), .Q(
        \register[2][28] ), .QN(n2393) );
  DFFRX1 \register_reg[2][27]  ( .D(n141), .CK(clk), .RN(n2253), .Q(
        \register[2][27] ), .QN(n2392) );
  DFFRX1 \register_reg[2][26]  ( .D(n140), .CK(clk), .RN(n2253), .Q(
        \register[2][26] ), .QN(n2391) );
  DFFRX1 \register_reg[2][25]  ( .D(n139), .CK(clk), .RN(n2253), .Q(
        \register[2][25] ), .QN(n2390) );
  DFFRX1 \register_reg[2][24]  ( .D(n138), .CK(clk), .RN(n2253), .Q(
        \register[2][24] ), .QN(n2389) );
  DFFRX1 \register_reg[2][23]  ( .D(n137), .CK(clk), .RN(n2253), .Q(
        \register[2][23] ), .QN(n2388) );
  DFFRX1 \register_reg[2][22]  ( .D(n136), .CK(clk), .RN(n2253), .Q(
        \register[2][22] ), .QN(n2387) );
  DFFRX1 \register_reg[2][21]  ( .D(n135), .CK(clk), .RN(n2253), .Q(
        \register[2][21] ), .QN(n2386) );
  DFFRX1 \register_reg[2][20]  ( .D(n134), .CK(clk), .RN(n2253), .Q(
        \register[2][20] ), .QN(n2385) );
  DFFRX1 \register_reg[2][19]  ( .D(n133), .CK(clk), .RN(n2253), .Q(
        \register[2][19] ), .QN(n2384) );
  DFFRX1 \register_reg[2][18]  ( .D(n132), .CK(clk), .RN(n2253), .Q(
        \register[2][18] ), .QN(n2383) );
  DFFRX1 \register_reg[2][17]  ( .D(n131), .CK(clk), .RN(n2253), .Q(
        \register[2][17] ), .QN(n2382) );
  DFFRX1 \register_reg[2][16]  ( .D(n130), .CK(clk), .RN(n2253), .Q(
        \register[2][16] ), .QN(n2381) );
  DFFRX1 \register_reg[2][15]  ( .D(n129), .CK(clk), .RN(n2253), .Q(
        \register[2][15] ), .QN(n2380) );
  DFFRX1 \register_reg[2][14]  ( .D(n128), .CK(clk), .RN(n2253), .Q(
        \register[2][14] ), .QN(n2379) );
  DFFRX1 \register_reg[2][13]  ( .D(n127), .CK(clk), .RN(n2253), .Q(
        \register[2][13] ), .QN(n2378) );
  DFFRX1 \register_reg[2][12]  ( .D(n126), .CK(clk), .RN(n2253), .Q(
        \register[2][12] ), .QN(n2377) );
  DFFRX1 \register_reg[2][11]  ( .D(n125), .CK(clk), .RN(n2253), .Q(
        \register[2][11] ), .QN(n2376) );
  DFFRX1 \register_reg[2][10]  ( .D(n124), .CK(clk), .RN(n2253), .Q(
        \register[2][10] ), .QN(n2375) );
  DFFRX1 \register_reg[2][9]  ( .D(n123), .CK(clk), .RN(n2253), .Q(
        \register[2][9] ), .QN(n2374) );
  DFFRX1 \register_reg[2][8]  ( .D(n122), .CK(clk), .RN(n2253), .Q(
        \register[2][8] ), .QN(n2373) );
  DFFRX1 \register_reg[2][7]  ( .D(n121), .CK(clk), .RN(n2253), .Q(
        \register[2][7] ), .QN(n2372) );
  DFFRX1 \register_reg[2][6]  ( .D(n120), .CK(clk), .RN(n2253), .Q(
        \register[2][6] ), .QN(n2371) );
  DFFRX1 \register_reg[2][5]  ( .D(n119), .CK(clk), .RN(n2253), .Q(
        \register[2][5] ), .QN(n2370) );
  DFFRX1 \register_reg[2][4]  ( .D(n118), .CK(clk), .RN(n2253), .Q(
        \register[2][4] ), .QN(n2369) );
  DFFRX1 \register_reg[2][3]  ( .D(n117), .CK(clk), .RN(n2253), .Q(
        \register[2][3] ), .QN(n2368) );
  DFFRX1 \register_reg[2][2]  ( .D(n116), .CK(clk), .RN(n2253), .Q(
        \register[2][2] ), .QN(n2367) );
  DFFRX1 \register_reg[2][1]  ( .D(n115), .CK(clk), .RN(n2253), .Q(
        \register[2][1] ), .QN(n2366) );
  DFFRX1 \register_reg[2][0]  ( .D(n114), .CK(clk), .RN(n2253), .Q(
        \register[2][0] ), .QN(n2365) );
  DFFRX1 \register_reg[1][1]  ( .D(n83), .CK(clk), .RN(n2253), .Q(
        \register[1][1] ), .QN(n2) );
  OAI22X1 U2 ( .A0(n1993), .A1(n2022), .B0(n1988), .B1(\register[1][0] ), .Y(
        n1951) );
  NOR3BXL U3 ( .AN(n53), .B(WriteReg[3]), .C(WriteReg[4]), .Y(n40) );
  NOR3BXL U4 ( .AN(n53), .B(WriteReg[4]), .C(n2431), .Y(n56) );
  MXI2X1 U5 ( .A(n3), .B(n4), .S0(n1455), .Y(ReadData1[0]) );
  MX4X1 U6 ( .A(n1607), .B(n1605), .C(n1606), .D(n1604), .S0(n1957), .S1(n1966), .Y(n1536) );
  MXI2X1 U7 ( .A(n1536), .B(n1537), .S0(n1952), .Y(ReadData2[0]) );
  MX4X1 U8 ( .A(n1603), .B(n1601), .C(n1602), .D(n1600), .S0(n1957), .S1(n1966), .Y(n1537) );
  OAI2BB2XL U9 ( .B0(n1993), .B1(n2021), .A0N(n1), .A1N(n2), .Y(n1948) );
  CLKINVX1 U10 ( .A(n1989), .Y(n1) );
  MXI2X1 U11 ( .A(n13), .B(n14), .S0(n1455), .Y(ReadData1[5]) );
  MXI4XL U12 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1519), .S1(n1488), .Y(
        n1139) );
  MXI4XL U13 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1517), .S1(n1488), .Y(
        n1107) );
  MXI4XL U14 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1518), .S1(n1488), .Y(
        n1115) );
  MXI4XL U15 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1518), .S1(n1488), .Y(
        n1123) );
  MXI4XL U16 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1519), .S1(n1488), .Y(
        n1131) );
  MXI4XL U17 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1519), .S1(n1488), .Y(
        n1147) );
  MXI4XL U18 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1519), .S1(n1488), .Y(
        n1138) );
  MXI4XL U19 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1517), .S1(n1488), .Y(
        n1106) );
  MXI4XL U20 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1518), .S1(n1488), .Y(
        n1114) );
  MXI4XL U21 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1518), .S1(n1488), .Y(
        n1122) );
  MXI4XL U22 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1518), .S1(n1488), .Y(
        n1130) );
  MXI4XL U23 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1519), .S1(n1488), .Y(
        n1146) );
  MXI4XL U24 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1520), .S1(n1489), .Y(
        n1155) );
  MXI4XL U25 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1517), .S1(n1487), .Y(
        n1105) );
  MXI4XL U26 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(\register[6][4] ), .D(\register[7][4] ), .S0(n1519), .S1(n1488), .Y(n1141) );
  MXI4XL U27 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1519), .S1(n1488), .Y(
        n1137) );
  MXI4XL U28 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(\register[6][0] ), .D(\register[7][0] ), .S0(n1517), .S1(n1488), .Y(n1109) );
  MXI4XL U29 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(\register[6][1] ), .D(\register[7][1] ), .S0(n1518), .S1(n1488), .Y(n1117) );
  MXI4XL U30 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1518), .S1(n1488), .Y(
        n1113) );
  MXI4XL U31 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(\register[6][2] ), .D(\register[7][2] ), .S0(n1518), .S1(n1488), .Y(n1125) );
  MXI4XL U32 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1518), .S1(n1488), .Y(
        n1121) );
  MXI4XL U33 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(\register[6][3] ), .D(\register[7][3] ), .S0(n1519), .S1(n1488), .Y(n1133) );
  MXI4XL U34 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1518), .S1(n1488), .Y(
        n1129) );
  MXI4XL U35 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1519), .S1(n1488), .Y(
        n1145) );
  MXI4XL U36 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1520), .S1(n1489), .Y(
        n1154) );
  MXI4XL U37 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(\register[6][6] ), .D(\register[7][6] ), .S0(n1520), .S1(n1489), .Y(n1157) );
  MXI4XL U38 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1520), .S1(n1489), .Y(
        n1153) );
  MXI4XL U39 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(\register[6][5] ), .D(\register[7][5] ), .S0(n1519), .S1(n1489), .Y(n1149) );
  MXI4XL U40 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1517), .S1(n1487), .Y(
        n1104) );
  MXI4XL U41 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1519), .S1(n1488), .Y(
        n1140) );
  MXI4XL U42 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1519), .S1(n1488), .Y(
        n1136) );
  MXI4XL U43 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1517), .S1(n1488), .Y(
        n1108) );
  MXI4XL U44 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1518), .S1(n1488), .Y(
        n1116) );
  MXI4XL U45 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1518), .S1(n1488), .Y(
        n1112) );
  MXI4XL U46 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1518), .S1(n1488), .Y(
        n1124) );
  MXI4XL U47 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1518), .S1(n1488), .Y(
        n1120) );
  MXI4XL U48 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1519), .S1(n1488), .Y(
        n1132) );
  MXI4XL U49 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1518), .S1(n1488), .Y(
        n1128) );
  MXI4XL U50 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1519), .S1(n1488), .Y(
        n1144) );
  MXI4XL U51 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1520), .S1(n1489), .Y(
        n1156) );
  MXI4XL U52 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1520), .S1(n1489), .Y(
        n1152) );
  MXI4XL U53 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1519), .S1(n1489), .Y(
        n1148) );
  NAND2X1 U54 ( .A(n52), .B(n40), .Y(n51) );
  NAND2X1 U55 ( .A(n56), .B(n52), .Y(n63) );
  NAND2X1 U56 ( .A(n65), .B(n52), .Y(n72) );
  NAND2X1 U57 ( .A(n74), .B(n52), .Y(n81) );
  NAND2X1 U58 ( .A(n39), .B(n40), .Y(n38) );
  NAND2X1 U59 ( .A(n42), .B(n40), .Y(n41) );
  NAND2X1 U60 ( .A(n44), .B(n40), .Y(n43) );
  NAND2X1 U61 ( .A(n46), .B(n40), .Y(n45) );
  NAND2X1 U62 ( .A(n48), .B(n40), .Y(n47) );
  NAND2X1 U63 ( .A(n50), .B(n40), .Y(n49) );
  NAND2X1 U64 ( .A(n56), .B(n39), .Y(n57) );
  NAND2X1 U65 ( .A(n56), .B(n42), .Y(n58) );
  NAND2X1 U66 ( .A(n56), .B(n44), .Y(n59) );
  NAND2X1 U67 ( .A(n56), .B(n46), .Y(n60) );
  NAND2X1 U68 ( .A(n56), .B(n48), .Y(n61) );
  NAND2X1 U69 ( .A(n56), .B(n50), .Y(n62) );
  NAND2X1 U70 ( .A(n55), .B(n56), .Y(n54) );
  NAND2X1 U71 ( .A(n65), .B(n46), .Y(n69) );
  NAND2X1 U72 ( .A(n65), .B(n48), .Y(n70) );
  NAND2X1 U73 ( .A(n65), .B(n50), .Y(n71) );
  NAND2X1 U74 ( .A(n74), .B(n46), .Y(n78) );
  NAND2X1 U75 ( .A(n74), .B(n48), .Y(n79) );
  NAND2X1 U76 ( .A(n74), .B(n50), .Y(n80) );
  NAND2X1 U77 ( .A(n65), .B(n42), .Y(n67) );
  NAND2X1 U78 ( .A(n65), .B(n44), .Y(n68) );
  NAND2X1 U79 ( .A(n74), .B(n42), .Y(n76) );
  NAND2X1 U80 ( .A(n74), .B(n44), .Y(n77) );
  NAND2X1 U81 ( .A(n65), .B(n39), .Y(n66) );
  NAND2X1 U82 ( .A(n74), .B(n39), .Y(n75) );
  NAND2X1 U83 ( .A(n65), .B(n55), .Y(n64) );
  NAND2X1 U84 ( .A(n74), .B(n55), .Y(n73) );
  NOR3X1 U85 ( .A(WriteReg[1]), .B(WriteReg[2]), .C(n2428), .Y(n39) );
  NOR3X1 U86 ( .A(WriteReg[0]), .B(WriteReg[2]), .C(n2429), .Y(n42) );
  NOR3X1 U87 ( .A(n2428), .B(WriteReg[2]), .C(n2429), .Y(n44) );
  NOR3X1 U88 ( .A(WriteReg[0]), .B(WriteReg[1]), .C(n2430), .Y(n46) );
  NOR3X1 U89 ( .A(n2428), .B(WriteReg[1]), .C(n2430), .Y(n48) );
  NOR3X1 U90 ( .A(n2429), .B(WriteReg[0]), .C(n2430), .Y(n50) );
  NOR3X1 U91 ( .A(WriteReg[1]), .B(WriteReg[2]), .C(WriteReg[0]), .Y(n55) );
  CLKINVX1 U92 ( .A(WriteReg[2]), .Y(n2430) );
  CLKINVX1 U93 ( .A(WriteReg[1]), .Y(n2429) );
  CLKINVX1 U94 ( .A(WriteReg[0]), .Y(n2428) );
  MXI4XL U95 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1517), .S1(n1487), .Y(
        n1103) );
  NOR2BXL U96 ( .AN(n1490), .B(\register[3][0] ), .Y(n1452) );
  MXI4XL U97 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1521), .S1(n1490), .Y(
        n1175) );
  MXI4XL U98 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1518), .S1(n1488), .Y(
        n1127) );
  MXI4XL U99 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1191) );
  MXI4XL U100 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1522), .S1(n1490), 
        .Y(n1207) );
  MXI4XL U101 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1518), .S1(n1488), .Y(
        n1119) );
  MXI4XL U102 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1521), .S1(n1490), 
        .Y(n1183) );
  MXI4XL U103 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1199) );
  MXI2X1 U104 ( .A(n5), .B(n6), .S0(n1455), .Y(ReadData1[1]) );
  MXI4XL U105 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1517), .S1(n1488), .Y(
        n1111) );
  MXI2X1 U106 ( .A(n31), .B(n32), .S0(n1456), .Y(ReadData1[14]) );
  MXI4XL U107 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1215) );
  MXI2X1 U108 ( .A(n35), .B(n36), .S0(n1456), .Y(ReadData1[16]) );
  MXI4XL U109 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1511), .S1(n1484), 
        .Y(n1231) );
  MXI2X1 U110 ( .A(n37), .B(n1074), .S0(n1456), .Y(ReadData1[17]) );
  MXI2X1 U111 ( .A(n1083), .B(n1084), .S0(n1457), .Y(ReadData1[22]) );
  MXI2X1 U112 ( .A(n1087), .B(n1088), .S0(n1457), .Y(ReadData1[24]) );
  MXI2X1 U113 ( .A(n1089), .B(n1090), .S0(n1457), .Y(ReadData1[25]) );
  MXI2X1 U114 ( .A(n11), .B(n12), .S0(n1455), .Y(ReadData1[4]) );
  MXI4XL U115 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1519), .S1(n1488), .Y(
        n1135) );
  MXI4XL U116 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1519), .S1(n1488), .Y(
        n1143) );
  MXI2X1 U117 ( .A(n15), .B(n16), .S0(n1455), .Y(ReadData1[6]) );
  MXI4XL U118 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1520), .S1(n1489), .Y(
        n1151) );
  MXI2X1 U119 ( .A(n17), .B(n18), .S0(n1455), .Y(ReadData1[7]) );
  MXI4XL U120 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1520), .S1(n1489), .Y(
        n1159) );
  NOR2BXL U121 ( .AN(n1491), .B(\register[3][1] ), .Y(n1449) );
  MXI2XL U122 ( .A(n2367), .B(n1446), .S0(n1528), .Y(n1447) );
  NOR2BXL U123 ( .AN(n1491), .B(\register[3][2] ), .Y(n1446) );
  MXI2XL U124 ( .A(n2368), .B(n1443), .S0(n1528), .Y(n1444) );
  NOR2BXL U125 ( .AN(n1491), .B(\register[3][3] ), .Y(n1443) );
  NOR2BXL U126 ( .AN(n1491), .B(\register[3][4] ), .Y(n1440) );
  NOR2BXL U127 ( .AN(n1491), .B(\register[3][5] ), .Y(n1437) );
  NOR2BXL U128 ( .AN(n1491), .B(\register[3][6] ), .Y(n1434) );
  MXI2XL U129 ( .A(n2373), .B(n1428), .S0(n1528), .Y(n1429) );
  NOR2BXL U130 ( .AN(n1491), .B(\register[3][8] ), .Y(n1428) );
  NOR2BXL U131 ( .AN(n1491), .B(\register[3][7] ), .Y(n1431) );
  MXI2XL U132 ( .A(n2374), .B(n1425), .S0(n1527), .Y(n1426) );
  NOR2BXL U133 ( .AN(n1491), .B(\register[3][9] ), .Y(n1425) );
  MXI2XL U134 ( .A(n2375), .B(n1422), .S0(n1527), .Y(n1423) );
  NOR2BXL U135 ( .AN(n1491), .B(\register[3][10] ), .Y(n1422) );
  MXI2XL U136 ( .A(n2376), .B(n1419), .S0(n1527), .Y(n1420) );
  NOR2BXL U137 ( .AN(n1491), .B(\register[3][11] ), .Y(n1419) );
  MXI2XL U138 ( .A(n2377), .B(n1416), .S0(n1527), .Y(n1417) );
  NOR2BXL U139 ( .AN(n1491), .B(\register[3][12] ), .Y(n1416) );
  MXI2XL U140 ( .A(n2378), .B(n1413), .S0(n1527), .Y(n1414) );
  NOR2BXL U141 ( .AN(n1491), .B(\register[3][13] ), .Y(n1413) );
  NOR2BXL U142 ( .AN(n1491), .B(\register[3][14] ), .Y(n1410) );
  MXI4XL U143 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1520), .S1(n1490), .Y(
        n1167) );
  MXI4XL U144 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1520), .S1(n1489), .Y(
        n1163) );
  MXI4XL U145 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1523), .S1(n1489), 
        .Y(n1211) );
  MXI4XL U146 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1219) );
  MXI4XL U147 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1511), .S1(n1485), 
        .Y(n1235) );
  MXI4XL U148 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1521), .S1(n1490), .Y(
        n1171) );
  MXI4XL U149 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1521), .S1(n1490), .Y(
        n1179) );
  MXI4XL U150 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1521), .S1(n1490), 
        .Y(n1187) );
  MXI4XL U151 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1195) );
  MXI4XL U152 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1203) );
  MXI4XL U153 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1520), .S1(n1489), .Y(
        n1162) );
  MXI4XL U154 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1523), .S1(n1489), 
        .Y(n1210) );
  MXI4XL U155 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1218) );
  MXI4XL U156 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1511), .S1(n1485), 
        .Y(n1234) );
  MXI4XL U157 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1521), .S1(n1490), .Y(
        n1170) );
  MXI4XL U158 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1521), .S1(n1490), .Y(
        n1178) );
  MXI4XL U159 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1521), .S1(n1490), 
        .Y(n1186) );
  MXI4XL U160 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1194) );
  MXI4XL U161 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1202) );
  MXI4XL U162 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1520), .S1(n1489), .Y(
        n1161) );
  MXI4XL U163 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1520), .S1(n1489), .Y(
        n1165) );
  MXI4XL U164 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1523), .S1(n1489), .Y(
        n1213) );
  MXI4XL U165 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1523), .S1(n1489), 
        .Y(n1209) );
  MXI4XL U166 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1217) );
  MXI4XL U167 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1523), .S1(n1489), .Y(
        n1221) );
  MXI4XL U168 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1511), .S1(n1485), .Y(
        n1237) );
  MXI4XL U169 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1521), .S1(n1490), .Y(
        n1173) );
  MXI4XL U170 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1521), .S1(n1490), .Y(
        n1169) );
  MXI4XL U171 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1521), .S1(n1490), .Y(
        n1181) );
  MXI4XL U172 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1521), .S1(n1490), .Y(
        n1177) );
  MXI4XL U173 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1522), .S1(n1490), .Y(
        n1189) );
  MXI4XL U174 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1521), .S1(n1490), 
        .Y(n1185) );
  MXI4XL U175 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1522), .S1(n1490), .Y(
        n1197) );
  MXI4XL U176 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1193) );
  MXI4XL U177 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1522), .S1(n1490), .Y(
        n1205) );
  MXI4XL U178 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1201) );
  MXI4XL U179 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1520), .S1(n1489), .Y(
        n1160) );
  MXI4XL U180 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1520), .S1(n1489), .Y(
        n1164) );
  MXI4XL U181 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1523), .S1(n1489), 
        .Y(n1212) );
  MXI4XL U182 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1523), .S1(n1489), 
        .Y(n1208) );
  MXI4XL U183 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1216) );
  MXI4XL U184 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1523), .S1(n1489), 
        .Y(n1220) );
  MXI4XL U185 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1511), .S1(n1485), 
        .Y(n1236) );
  MXI4XL U186 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1521), .S1(n1490), .Y(
        n1172) );
  MXI4XL U187 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1520), .S1(n1490), .Y(
        n1168) );
  MXI4XL U188 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1521), .S1(n1490), .Y(
        n1180) );
  MXI4XL U189 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1521), .S1(n1490), .Y(
        n1176) );
  MXI4XL U190 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1522), .S1(n1490), 
        .Y(n1188) );
  MXI4XL U191 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1521), .S1(n1490), 
        .Y(n1184) );
  MXI4XL U192 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1196) );
  MXI4XL U193 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1522), .S1(n1490), 
        .Y(n1192) );
  MXI4XL U194 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1204) );
  MXI4XL U195 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1522), .S1(n1490), 
        .Y(n1200) );
  MXI4XL U196 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1511), .S1(n1484), 
        .Y(n1233) );
  MXI4XL U197 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1511), .S1(n1484), 
        .Y(n1232) );
  MXI2X1 U198 ( .A(n1099), .B(n1100), .S0(n1457), .Y(ReadData1[30]) );
  CLKINVX1 U199 ( .A(n2350), .Y(n2254) );
  CLKINVX1 U200 ( .A(n2350), .Y(n2255) );
  CLKINVX1 U201 ( .A(n2349), .Y(n2256) );
  CLKINVX1 U202 ( .A(n2349), .Y(n2257) );
  CLKINVX1 U203 ( .A(n2349), .Y(n2258) );
  CLKINVX1 U204 ( .A(n2348), .Y(n2259) );
  CLKINVX1 U205 ( .A(n2348), .Y(n2260) );
  CLKINVX1 U206 ( .A(n2348), .Y(n2261) );
  CLKINVX1 U207 ( .A(n2347), .Y(n2262) );
  CLKINVX1 U208 ( .A(n2347), .Y(n2263) );
  CLKINVX1 U209 ( .A(n2347), .Y(n2264) );
  CLKINVX1 U210 ( .A(n2346), .Y(n2265) );
  CLKINVX1 U211 ( .A(n2346), .Y(n2266) );
  CLKINVX1 U212 ( .A(n2346), .Y(n2267) );
  CLKINVX1 U213 ( .A(n2345), .Y(n2268) );
  CLKINVX1 U214 ( .A(n2345), .Y(n2269) );
  CLKINVX1 U215 ( .A(n2345), .Y(n2270) );
  CLKINVX1 U216 ( .A(n2344), .Y(n2271) );
  CLKINVX1 U217 ( .A(n2344), .Y(n2272) );
  CLKINVX1 U218 ( .A(n2344), .Y(n2273) );
  CLKINVX1 U219 ( .A(n2343), .Y(n2274) );
  CLKINVX1 U220 ( .A(n2343), .Y(n2275) );
  CLKINVX1 U221 ( .A(n2343), .Y(n2276) );
  CLKINVX1 U222 ( .A(n2342), .Y(n2277) );
  CLKINVX1 U223 ( .A(n2342), .Y(n2278) );
  CLKINVX1 U224 ( .A(n2342), .Y(n2279) );
  CLKINVX1 U225 ( .A(n2341), .Y(n2280) );
  CLKINVX1 U226 ( .A(n2341), .Y(n2281) );
  CLKINVX1 U227 ( .A(n2341), .Y(n2282) );
  CLKINVX1 U228 ( .A(n2340), .Y(n2283) );
  CLKINVX1 U229 ( .A(n2340), .Y(n2284) );
  CLKINVX1 U230 ( .A(n2340), .Y(n2285) );
  CLKINVX1 U231 ( .A(n2339), .Y(n2286) );
  CLKINVX1 U232 ( .A(n2339), .Y(n2287) );
  CLKINVX1 U233 ( .A(n2339), .Y(n2288) );
  CLKINVX1 U234 ( .A(n2338), .Y(n2289) );
  CLKINVX1 U235 ( .A(n2338), .Y(n2290) );
  CLKINVX1 U236 ( .A(n2338), .Y(n2291) );
  CLKINVX1 U237 ( .A(n2337), .Y(n2292) );
  CLKINVX1 U238 ( .A(n2337), .Y(n2293) );
  CLKINVX1 U239 ( .A(n2337), .Y(n2294) );
  CLKINVX1 U240 ( .A(n2336), .Y(n2295) );
  CLKINVX1 U241 ( .A(n2336), .Y(n2296) );
  CLKINVX1 U242 ( .A(n2336), .Y(n2297) );
  CLKINVX1 U243 ( .A(n2335), .Y(n2298) );
  CLKINVX1 U244 ( .A(n2335), .Y(n2299) );
  CLKINVX1 U245 ( .A(n2335), .Y(n2300) );
  CLKINVX1 U246 ( .A(n2334), .Y(n2301) );
  CLKINVX1 U247 ( .A(n2334), .Y(n2302) );
  CLKINVX1 U248 ( .A(n2334), .Y(n2303) );
  CLKINVX1 U249 ( .A(n2333), .Y(n2304) );
  CLKINVX1 U250 ( .A(n2333), .Y(n2305) );
  CLKINVX1 U251 ( .A(n2333), .Y(n2306) );
  CLKINVX1 U252 ( .A(n2332), .Y(n2307) );
  CLKINVX1 U253 ( .A(n2332), .Y(n2308) );
  CLKINVX1 U254 ( .A(n2332), .Y(n2309) );
  CLKINVX1 U255 ( .A(n2331), .Y(n2310) );
  CLKINVX1 U256 ( .A(n2331), .Y(n2311) );
  CLKINVX1 U257 ( .A(n2331), .Y(n2312) );
  CLKINVX1 U258 ( .A(n2330), .Y(n2313) );
  CLKINVX1 U259 ( .A(n2330), .Y(n2314) );
  CLKINVX1 U260 ( .A(n2330), .Y(n2315) );
  CLKINVX1 U261 ( .A(n2329), .Y(n2316) );
  CLKINVX1 U262 ( .A(n2329), .Y(n2317) );
  CLKINVX1 U263 ( .A(n2329), .Y(n2318) );
  CLKINVX1 U264 ( .A(n2328), .Y(n2319) );
  CLKINVX1 U265 ( .A(n2328), .Y(n2320) );
  CLKINVX1 U266 ( .A(n2328), .Y(n2321) );
  CLKINVX1 U267 ( .A(n2327), .Y(n2322) );
  CLKINVX1 U268 ( .A(n2327), .Y(n2323) );
  CLKINVX1 U269 ( .A(n2327), .Y(n2324) );
  CLKINVX1 U270 ( .A(n2326), .Y(n2325) );
  CLKBUFX3 U271 ( .A(n1503), .Y(n1525) );
  CLKBUFX3 U272 ( .A(n2000), .Y(n2022) );
  CLKBUFX3 U273 ( .A(n1506), .Y(n1519) );
  CLKBUFX3 U274 ( .A(n1506), .Y(n1520) );
  CLKBUFX3 U275 ( .A(n1505), .Y(n1521) );
  CLKBUFX3 U276 ( .A(n1505), .Y(n1522) );
  CLKBUFX3 U277 ( .A(n1504), .Y(n1523) );
  CLKBUFX3 U278 ( .A(n1510), .Y(n1511) );
  CLKBUFX3 U279 ( .A(n1510), .Y(n1512) );
  CLKBUFX3 U280 ( .A(n1509), .Y(n1513) );
  CLKBUFX3 U281 ( .A(n1509), .Y(n1514) );
  CLKBUFX3 U282 ( .A(n1508), .Y(n1515) );
  CLKBUFX3 U283 ( .A(n1507), .Y(n1518) );
  CLKBUFX3 U284 ( .A(n1508), .Y(n1516) );
  CLKBUFX3 U285 ( .A(n1507), .Y(n1517) );
  CLKBUFX3 U286 ( .A(n2004), .Y(n2015) );
  CLKBUFX3 U287 ( .A(n2003), .Y(n2016) );
  CLKBUFX3 U288 ( .A(n2002), .Y(n2018) );
  CLKBUFX3 U289 ( .A(n2002), .Y(n2019) );
  CLKBUFX3 U290 ( .A(n2003), .Y(n2017) );
  CLKBUFX3 U291 ( .A(n2001), .Y(n2020) );
  CLKBUFX3 U292 ( .A(n2007), .Y(n2008) );
  CLKBUFX3 U293 ( .A(n2007), .Y(n2009) );
  CLKBUFX3 U294 ( .A(n2006), .Y(n2010) );
  CLKBUFX3 U295 ( .A(n2005), .Y(n2012) );
  CLKBUFX3 U296 ( .A(n2005), .Y(n2013) );
  CLKBUFX3 U297 ( .A(n2006), .Y(n2011) );
  CLKBUFX3 U298 ( .A(n2004), .Y(n2014) );
  CLKBUFX3 U299 ( .A(n1504), .Y(n1524) );
  CLKBUFX3 U300 ( .A(n2001), .Y(n2021) );
  CLKBUFX3 U301 ( .A(n1503), .Y(n1526) );
  CLKBUFX3 U302 ( .A(n2000), .Y(n2023) );
  CLKBUFX3 U303 ( .A(n1478), .Y(n1494) );
  CLKBUFX3 U304 ( .A(n1975), .Y(n1991) );
  CLKBUFX3 U305 ( .A(n1479), .Y(n1493) );
  CLKBUFX3 U306 ( .A(n1479), .Y(n1492) );
  CLKBUFX3 U307 ( .A(n1976), .Y(n1989) );
  CLKBUFX3 U308 ( .A(n1976), .Y(n1990) );
  CLKBUFX3 U309 ( .A(n1480), .Y(n1490) );
  CLKBUFX3 U310 ( .A(n1977), .Y(n1987) );
  CLKBUFX3 U311 ( .A(n1481), .Y(n1489) );
  CLKBUFX3 U312 ( .A(n1483), .Y(n1485) );
  CLKBUFX3 U313 ( .A(n1482), .Y(n1486) );
  CLKBUFX3 U314 ( .A(n1481), .Y(n1488) );
  CLKBUFX3 U315 ( .A(n1482), .Y(n1487) );
  CLKBUFX3 U316 ( .A(n1978), .Y(n1985) );
  CLKBUFX3 U317 ( .A(n1980), .Y(n1982) );
  CLKBUFX3 U318 ( .A(n1979), .Y(n1983) );
  CLKBUFX3 U319 ( .A(n1978), .Y(n1986) );
  CLKBUFX3 U320 ( .A(n1979), .Y(n1984) );
  CLKBUFX3 U321 ( .A(n1480), .Y(n1491) );
  CLKBUFX3 U322 ( .A(n1977), .Y(n1988) );
  CLKBUFX3 U323 ( .A(n1478), .Y(n1495) );
  CLKBUFX3 U324 ( .A(n1975), .Y(n1992) );
  CLKBUFX3 U325 ( .A(n2352), .Y(n2349) );
  CLKBUFX3 U326 ( .A(n2352), .Y(n2348) );
  CLKBUFX3 U327 ( .A(n2353), .Y(n2347) );
  CLKBUFX3 U328 ( .A(n2353), .Y(n2346) );
  CLKBUFX3 U329 ( .A(n2354), .Y(n2345) );
  CLKBUFX3 U330 ( .A(n2354), .Y(n2344) );
  CLKBUFX3 U331 ( .A(n2355), .Y(n2343) );
  CLKBUFX3 U332 ( .A(n2355), .Y(n2342) );
  CLKBUFX3 U333 ( .A(n2356), .Y(n2341) );
  CLKBUFX3 U334 ( .A(n2356), .Y(n2340) );
  CLKBUFX3 U335 ( .A(n2357), .Y(n2339) );
  CLKBUFX3 U336 ( .A(n2357), .Y(n2338) );
  CLKBUFX3 U337 ( .A(n2358), .Y(n2337) );
  CLKBUFX3 U338 ( .A(n2358), .Y(n2336) );
  CLKBUFX3 U339 ( .A(n2359), .Y(n2335) );
  CLKBUFX3 U340 ( .A(n2359), .Y(n2334) );
  CLKBUFX3 U341 ( .A(n2360), .Y(n2333) );
  CLKBUFX3 U342 ( .A(n2360), .Y(n2332) );
  CLKBUFX3 U343 ( .A(n2361), .Y(n2331) );
  CLKBUFX3 U344 ( .A(n2361), .Y(n2330) );
  CLKBUFX3 U345 ( .A(n2362), .Y(n2329) );
  CLKBUFX3 U346 ( .A(n2362), .Y(n2328) );
  CLKBUFX3 U347 ( .A(n2363), .Y(n2327) );
  CLKBUFX3 U348 ( .A(n2363), .Y(n2326) );
  CLKBUFX3 U349 ( .A(n2351), .Y(n2350) );
  CLKBUFX3 U350 ( .A(n1483), .Y(n1484) );
  CLKBUFX3 U351 ( .A(n1980), .Y(n1981) );
  CLKBUFX3 U352 ( .A(n38), .Y(n2251) );
  CLKBUFX3 U353 ( .A(n1502), .Y(n1528) );
  CLKBUFX3 U354 ( .A(n1502), .Y(n1527) );
  CLKBUFX3 U355 ( .A(n1999), .Y(n2024) );
  CLKBUFX3 U356 ( .A(n1999), .Y(n2025) );
  CLKBUFX3 U357 ( .A(n38), .Y(n2250) );
  CLKBUFX3 U358 ( .A(n38), .Y(n2249) );
  CLKBUFX3 U359 ( .A(n57), .Y(n2219) );
  CLKBUFX3 U360 ( .A(n58), .Y(n2215) );
  CLKBUFX3 U361 ( .A(n59), .Y(n2211) );
  CLKBUFX3 U362 ( .A(n60), .Y(n2207) );
  CLKBUFX3 U363 ( .A(n61), .Y(n2203) );
  CLKBUFX3 U364 ( .A(n62), .Y(n2199) );
  CLKBUFX3 U365 ( .A(n63), .Y(n2195) );
  CLKBUFX3 U366 ( .A(n54), .Y(n2223) );
  CLKBUFX3 U367 ( .A(n57), .Y(n2218) );
  CLKBUFX3 U368 ( .A(n57), .Y(n2217) );
  CLKBUFX3 U369 ( .A(n58), .Y(n2214) );
  CLKBUFX3 U370 ( .A(n58), .Y(n2213) );
  CLKBUFX3 U371 ( .A(n59), .Y(n2210) );
  CLKBUFX3 U372 ( .A(n59), .Y(n2209) );
  CLKBUFX3 U373 ( .A(n60), .Y(n2206) );
  CLKBUFX3 U374 ( .A(n60), .Y(n2205) );
  CLKBUFX3 U375 ( .A(n61), .Y(n2202) );
  CLKBUFX3 U376 ( .A(n61), .Y(n2201) );
  CLKBUFX3 U377 ( .A(n62), .Y(n2198) );
  CLKBUFX3 U378 ( .A(n62), .Y(n2197) );
  CLKBUFX3 U379 ( .A(n63), .Y(n2194) );
  CLKBUFX3 U380 ( .A(n63), .Y(n2193) );
  CLKBUFX3 U381 ( .A(n41), .Y(n2247) );
  CLKBUFX3 U382 ( .A(n43), .Y(n2243) );
  CLKBUFX3 U383 ( .A(n45), .Y(n2239) );
  CLKBUFX3 U384 ( .A(n47), .Y(n2235) );
  CLKBUFX3 U385 ( .A(n49), .Y(n2231) );
  CLKBUFX3 U386 ( .A(n51), .Y(n2227) );
  CLKBUFX3 U387 ( .A(n54), .Y(n2222) );
  CLKBUFX3 U388 ( .A(n54), .Y(n2221) );
  CLKBUFX3 U389 ( .A(n66), .Y(n2187) );
  CLKBUFX3 U390 ( .A(n67), .Y(n2183) );
  CLKBUFX3 U391 ( .A(n68), .Y(n2179) );
  CLKBUFX3 U392 ( .A(n69), .Y(n2175) );
  CLKBUFX3 U393 ( .A(n70), .Y(n2171) );
  CLKBUFX3 U394 ( .A(n71), .Y(n2167) );
  CLKBUFX3 U395 ( .A(n72), .Y(n2163) );
  CLKBUFX3 U396 ( .A(n75), .Y(n2155) );
  CLKBUFX3 U397 ( .A(n76), .Y(n2151) );
  CLKBUFX3 U398 ( .A(n77), .Y(n2147) );
  CLKBUFX3 U399 ( .A(n78), .Y(n2143) );
  CLKBUFX3 U400 ( .A(n79), .Y(n2139) );
  CLKBUFX3 U401 ( .A(n80), .Y(n2135) );
  CLKBUFX3 U402 ( .A(n81), .Y(n2131) );
  CLKBUFX3 U403 ( .A(n64), .Y(n2191) );
  CLKBUFX3 U404 ( .A(n73), .Y(n2159) );
  CLKBUFX3 U405 ( .A(n41), .Y(n2246) );
  CLKBUFX3 U406 ( .A(n41), .Y(n2245) );
  CLKBUFX3 U407 ( .A(n43), .Y(n2242) );
  CLKBUFX3 U408 ( .A(n43), .Y(n2241) );
  CLKBUFX3 U409 ( .A(n45), .Y(n2238) );
  CLKBUFX3 U410 ( .A(n45), .Y(n2237) );
  CLKBUFX3 U411 ( .A(n47), .Y(n2234) );
  CLKBUFX3 U412 ( .A(n47), .Y(n2233) );
  CLKBUFX3 U413 ( .A(n49), .Y(n2230) );
  CLKBUFX3 U414 ( .A(n49), .Y(n2229) );
  CLKBUFX3 U415 ( .A(n51), .Y(n2226) );
  CLKBUFX3 U416 ( .A(n51), .Y(n2225) );
  CLKBUFX3 U417 ( .A(n66), .Y(n2186) );
  CLKBUFX3 U418 ( .A(n66), .Y(n2185) );
  CLKBUFX3 U419 ( .A(n67), .Y(n2182) );
  CLKBUFX3 U420 ( .A(n67), .Y(n2181) );
  CLKBUFX3 U421 ( .A(n68), .Y(n2178) );
  CLKBUFX3 U422 ( .A(n68), .Y(n2177) );
  CLKBUFX3 U423 ( .A(n69), .Y(n2174) );
  CLKBUFX3 U424 ( .A(n69), .Y(n2173) );
  CLKBUFX3 U425 ( .A(n70), .Y(n2170) );
  CLKBUFX3 U426 ( .A(n70), .Y(n2169) );
  CLKBUFX3 U427 ( .A(n71), .Y(n2166) );
  CLKBUFX3 U428 ( .A(n71), .Y(n2165) );
  CLKBUFX3 U429 ( .A(n72), .Y(n2162) );
  CLKBUFX3 U430 ( .A(n72), .Y(n2161) );
  CLKBUFX3 U431 ( .A(n75), .Y(n2154) );
  CLKBUFX3 U432 ( .A(n75), .Y(n2153) );
  CLKBUFX3 U433 ( .A(n76), .Y(n2150) );
  CLKBUFX3 U434 ( .A(n76), .Y(n2149) );
  CLKBUFX3 U435 ( .A(n77), .Y(n2146) );
  CLKBUFX3 U436 ( .A(n77), .Y(n2145) );
  CLKBUFX3 U437 ( .A(n78), .Y(n2142) );
  CLKBUFX3 U438 ( .A(n78), .Y(n2141) );
  CLKBUFX3 U439 ( .A(n79), .Y(n2138) );
  CLKBUFX3 U440 ( .A(n79), .Y(n2137) );
  CLKBUFX3 U441 ( .A(n80), .Y(n2134) );
  CLKBUFX3 U442 ( .A(n80), .Y(n2133) );
  CLKBUFX3 U443 ( .A(n81), .Y(n2130) );
  CLKBUFX3 U444 ( .A(n81), .Y(n2129) );
  CLKBUFX3 U445 ( .A(n64), .Y(n2190) );
  CLKBUFX3 U446 ( .A(n64), .Y(n2189) );
  CLKBUFX3 U447 ( .A(n73), .Y(n2158) );
  CLKBUFX3 U448 ( .A(n73), .Y(n2157) );
  CLKBUFX3 U449 ( .A(n57), .Y(n2220) );
  CLKBUFX3 U450 ( .A(n58), .Y(n2216) );
  CLKBUFX3 U451 ( .A(n59), .Y(n2212) );
  CLKBUFX3 U452 ( .A(n60), .Y(n2208) );
  CLKBUFX3 U453 ( .A(n61), .Y(n2204) );
  CLKBUFX3 U454 ( .A(n62), .Y(n2200) );
  CLKBUFX3 U455 ( .A(n63), .Y(n2196) );
  CLKBUFX3 U456 ( .A(n54), .Y(n2224) );
  CLKBUFX3 U457 ( .A(n41), .Y(n2248) );
  CLKBUFX3 U458 ( .A(n43), .Y(n2244) );
  CLKBUFX3 U459 ( .A(n45), .Y(n2240) );
  CLKBUFX3 U460 ( .A(n47), .Y(n2236) );
  CLKBUFX3 U461 ( .A(n49), .Y(n2232) );
  CLKBUFX3 U462 ( .A(n51), .Y(n2228) );
  CLKBUFX3 U463 ( .A(n66), .Y(n2188) );
  CLKBUFX3 U464 ( .A(n67), .Y(n2184) );
  CLKBUFX3 U465 ( .A(n68), .Y(n2180) );
  CLKBUFX3 U466 ( .A(n69), .Y(n2176) );
  CLKBUFX3 U467 ( .A(n70), .Y(n2172) );
  CLKBUFX3 U468 ( .A(n71), .Y(n2168) );
  CLKBUFX3 U469 ( .A(n72), .Y(n2164) );
  CLKBUFX3 U470 ( .A(n75), .Y(n2156) );
  CLKBUFX3 U471 ( .A(n76), .Y(n2152) );
  CLKBUFX3 U472 ( .A(n77), .Y(n2148) );
  CLKBUFX3 U473 ( .A(n78), .Y(n2144) );
  CLKBUFX3 U474 ( .A(n79), .Y(n2140) );
  CLKBUFX3 U475 ( .A(n80), .Y(n2136) );
  CLKBUFX3 U476 ( .A(n81), .Y(n2132) );
  CLKBUFX3 U477 ( .A(n64), .Y(n2192) );
  CLKBUFX3 U478 ( .A(n73), .Y(n2160) );
  CLKBUFX3 U479 ( .A(n38), .Y(n2252) );
  CLKBUFX3 U480 ( .A(n2357), .Y(n2351) );
  CLKBUFX3 U481 ( .A(n2358), .Y(n2352) );
  CLKBUFX3 U482 ( .A(n2359), .Y(n2353) );
  CLKBUFX3 U483 ( .A(n2360), .Y(n2354) );
  CLKBUFX3 U484 ( .A(n2361), .Y(n2355) );
  CLKBUFX3 U485 ( .A(n2362), .Y(n2356) );
  CLKBUFX3 U486 ( .A(n2364), .Y(n2357) );
  CLKBUFX3 U487 ( .A(n2364), .Y(n2358) );
  CLKBUFX3 U488 ( .A(n2364), .Y(n2359) );
  CLKBUFX3 U489 ( .A(n2364), .Y(n2360) );
  CLKBUFX3 U490 ( .A(n2364), .Y(n2361) );
  CLKBUFX3 U491 ( .A(n2364), .Y(n2362) );
  CLKBUFX3 U492 ( .A(n2364), .Y(n2363) );
  CLKBUFX3 U493 ( .A(n1533), .Y(n1506) );
  CLKBUFX3 U494 ( .A(n1533), .Y(n1505) );
  CLKBUFX3 U495 ( .A(n1532), .Y(n1504) );
  CLKBUFX3 U496 ( .A(n1500), .Y(n1481) );
  CLKBUFX3 U497 ( .A(n1501), .Y(n1483) );
  CLKBUFX3 U498 ( .A(n1535), .Y(n1510) );
  CLKBUFX3 U499 ( .A(n1535), .Y(n1509) );
  CLKBUFX3 U500 ( .A(n1499), .Y(n1478) );
  CLKBUFX3 U501 ( .A(n1501), .Y(n1482) );
  CLKBUFX3 U502 ( .A(n1534), .Y(n1508) );
  CLKBUFX3 U503 ( .A(n1499), .Y(n1479) );
  CLKBUFX3 U504 ( .A(n1532), .Y(n1503) );
  CLKBUFX3 U505 ( .A(n1534), .Y(n1507) );
  CLKBUFX3 U506 ( .A(n1500), .Y(n1480) );
  CLKBUFX3 U507 ( .A(n1997), .Y(n1977) );
  CLKBUFX3 U508 ( .A(n1996), .Y(n1976) );
  CLKBUFX3 U509 ( .A(n2029), .Y(n2000) );
  CLKBUFX3 U510 ( .A(n1996), .Y(n1975) );
  CLKBUFX3 U511 ( .A(n2030), .Y(n2002) );
  CLKBUFX3 U512 ( .A(n2030), .Y(n2003) );
  CLKBUFX3 U513 ( .A(n2032), .Y(n2007) );
  CLKBUFX3 U514 ( .A(n1998), .Y(n1980) );
  CLKBUFX3 U515 ( .A(n2031), .Y(n2005) );
  CLKBUFX3 U516 ( .A(n2032), .Y(n2006) );
  CLKBUFX3 U517 ( .A(n2029), .Y(n2001) );
  CLKBUFX3 U518 ( .A(n1997), .Y(n1978) );
  CLKBUFX3 U519 ( .A(n2031), .Y(n2004) );
  CLKBUFX3 U520 ( .A(n1998), .Y(n1979) );
  CLKBUFX3 U521 ( .A(n2432), .Y(n2127) );
  CLKBUFX3 U522 ( .A(n2427), .Y(n2124) );
  CLKBUFX3 U523 ( .A(n2426), .Y(n2121) );
  CLKBUFX3 U524 ( .A(n2425), .Y(n2118) );
  CLKBUFX3 U525 ( .A(n2424), .Y(n2115) );
  CLKBUFX3 U526 ( .A(n2423), .Y(n2112) );
  CLKBUFX3 U527 ( .A(n2422), .Y(n2109) );
  CLKBUFX3 U528 ( .A(n2421), .Y(n2106) );
  CLKBUFX3 U529 ( .A(n2420), .Y(n2103) );
  CLKBUFX3 U530 ( .A(n2419), .Y(n2100) );
  CLKBUFX3 U531 ( .A(n2418), .Y(n2097) );
  CLKBUFX3 U532 ( .A(n2417), .Y(n2094) );
  CLKBUFX3 U533 ( .A(n2416), .Y(n2091) );
  CLKBUFX3 U534 ( .A(n2415), .Y(n2088) );
  CLKBUFX3 U535 ( .A(n2414), .Y(n2085) );
  CLKBUFX3 U536 ( .A(n2413), .Y(n2082) );
  CLKBUFX3 U537 ( .A(n2412), .Y(n2079) );
  CLKBUFX3 U538 ( .A(n2411), .Y(n2076) );
  CLKBUFX3 U539 ( .A(n2410), .Y(n2073) );
  CLKBUFX3 U540 ( .A(n2409), .Y(n2070) );
  CLKBUFX3 U541 ( .A(n2408), .Y(n2067) );
  CLKBUFX3 U542 ( .A(n2407), .Y(n2064) );
  CLKBUFX3 U543 ( .A(n2406), .Y(n2061) );
  CLKBUFX3 U544 ( .A(n2405), .Y(n2058) );
  CLKBUFX3 U545 ( .A(n2404), .Y(n2055) );
  CLKBUFX3 U546 ( .A(n2403), .Y(n2052) );
  CLKBUFX3 U547 ( .A(n2402), .Y(n2049) );
  CLKBUFX3 U548 ( .A(n2401), .Y(n2046) );
  CLKBUFX3 U549 ( .A(n2400), .Y(n2043) );
  CLKBUFX3 U550 ( .A(n2399), .Y(n2040) );
  CLKBUFX3 U551 ( .A(n2398), .Y(n2037) );
  CLKBUFX3 U552 ( .A(n2397), .Y(n2034) );
  CLKBUFX3 U553 ( .A(n2432), .Y(n2126) );
  CLKBUFX3 U554 ( .A(n2427), .Y(n2123) );
  CLKBUFX3 U555 ( .A(n2426), .Y(n2120) );
  CLKBUFX3 U556 ( .A(n2425), .Y(n2117) );
  CLKBUFX3 U557 ( .A(n2424), .Y(n2114) );
  CLKBUFX3 U558 ( .A(n2423), .Y(n2111) );
  CLKBUFX3 U559 ( .A(n2422), .Y(n2108) );
  CLKBUFX3 U560 ( .A(n2421), .Y(n2105) );
  CLKBUFX3 U561 ( .A(n2420), .Y(n2102) );
  CLKBUFX3 U562 ( .A(n2419), .Y(n2099) );
  CLKBUFX3 U563 ( .A(n2418), .Y(n2096) );
  CLKBUFX3 U564 ( .A(n2417), .Y(n2093) );
  CLKBUFX3 U565 ( .A(n2416), .Y(n2090) );
  CLKBUFX3 U566 ( .A(n2415), .Y(n2087) );
  CLKBUFX3 U567 ( .A(n2414), .Y(n2084) );
  CLKBUFX3 U568 ( .A(n2413), .Y(n2081) );
  CLKBUFX3 U569 ( .A(n2412), .Y(n2078) );
  CLKBUFX3 U570 ( .A(n2411), .Y(n2075) );
  CLKBUFX3 U571 ( .A(n2410), .Y(n2072) );
  CLKBUFX3 U572 ( .A(n2409), .Y(n2069) );
  CLKBUFX3 U573 ( .A(n2408), .Y(n2066) );
  CLKBUFX3 U574 ( .A(n2407), .Y(n2063) );
  CLKBUFX3 U575 ( .A(n2406), .Y(n2060) );
  CLKBUFX3 U576 ( .A(n2405), .Y(n2057) );
  CLKBUFX3 U577 ( .A(n2404), .Y(n2054) );
  CLKBUFX3 U578 ( .A(n2403), .Y(n2051) );
  CLKBUFX3 U579 ( .A(n2402), .Y(n2048) );
  CLKBUFX3 U580 ( .A(n2401), .Y(n2045) );
  CLKBUFX3 U581 ( .A(n2400), .Y(n2042) );
  CLKBUFX3 U582 ( .A(n2399), .Y(n2039) );
  CLKBUFX3 U583 ( .A(n2398), .Y(n2036) );
  CLKBUFX3 U584 ( .A(n2397), .Y(n2033) );
  CLKBUFX3 U585 ( .A(n2432), .Y(n2128) );
  CLKBUFX3 U586 ( .A(n2427), .Y(n2125) );
  CLKBUFX3 U587 ( .A(n2426), .Y(n2122) );
  CLKBUFX3 U588 ( .A(n2425), .Y(n2119) );
  CLKBUFX3 U589 ( .A(n2424), .Y(n2116) );
  CLKBUFX3 U590 ( .A(n2423), .Y(n2113) );
  CLKBUFX3 U591 ( .A(n2422), .Y(n2110) );
  CLKBUFX3 U592 ( .A(n2421), .Y(n2107) );
  CLKBUFX3 U593 ( .A(n2420), .Y(n2104) );
  CLKBUFX3 U594 ( .A(n2419), .Y(n2101) );
  CLKBUFX3 U595 ( .A(n2418), .Y(n2098) );
  CLKBUFX3 U596 ( .A(n2417), .Y(n2095) );
  CLKBUFX3 U597 ( .A(n2416), .Y(n2092) );
  CLKBUFX3 U598 ( .A(n2415), .Y(n2089) );
  CLKBUFX3 U599 ( .A(n2414), .Y(n2086) );
  CLKBUFX3 U600 ( .A(n2413), .Y(n2083) );
  CLKBUFX3 U601 ( .A(n2412), .Y(n2080) );
  CLKBUFX3 U602 ( .A(n2411), .Y(n2077) );
  CLKBUFX3 U603 ( .A(n2410), .Y(n2074) );
  CLKBUFX3 U604 ( .A(n2409), .Y(n2071) );
  CLKBUFX3 U605 ( .A(n2408), .Y(n2068) );
  CLKBUFX3 U606 ( .A(n2407), .Y(n2065) );
  CLKBUFX3 U607 ( .A(n2406), .Y(n2062) );
  CLKBUFX3 U608 ( .A(n2405), .Y(n2059) );
  CLKBUFX3 U609 ( .A(n2404), .Y(n2056) );
  CLKBUFX3 U610 ( .A(n2403), .Y(n2053) );
  CLKBUFX3 U611 ( .A(n2402), .Y(n2050) );
  CLKBUFX3 U612 ( .A(n2401), .Y(n2047) );
  CLKBUFX3 U613 ( .A(n2400), .Y(n2044) );
  CLKBUFX3 U614 ( .A(n2399), .Y(n2041) );
  CLKBUFX3 U615 ( .A(n2398), .Y(n2038) );
  CLKBUFX3 U616 ( .A(n2397), .Y(n2035) );
  NOR3X1 U617 ( .A(n2429), .B(n2428), .C(n2430), .Y(n52) );
  CLKBUFX3 U618 ( .A(n1466), .Y(n1461) );
  CLKBUFX3 U619 ( .A(n1467), .Y(n1462) );
  CLKBUFX3 U620 ( .A(n1467), .Y(n1463) );
  CLKBUFX3 U621 ( .A(n1468), .Y(n1464) );
  CLKBUFX3 U622 ( .A(n1468), .Y(n1465) );
  CLKBUFX3 U623 ( .A(n1963), .Y(n1958) );
  CLKBUFX3 U624 ( .A(n1964), .Y(n1959) );
  CLKBUFX3 U625 ( .A(n1964), .Y(n1960) );
  CLKBUFX3 U626 ( .A(n1965), .Y(n1961) );
  CLKBUFX3 U627 ( .A(n1965), .Y(n1962) );
  CLKBUFX3 U628 ( .A(n1477), .Y(n1496) );
  CLKBUFX3 U629 ( .A(n1498), .Y(n1477) );
  CLKBUFX3 U630 ( .A(n1497), .Y(n1498) );
  CLKBUFX3 U631 ( .A(n1974), .Y(n1993) );
  CLKBUFX3 U632 ( .A(n1995), .Y(n1974) );
  CLKBUFX3 U633 ( .A(n1994), .Y(n1995) );
  CLKBUFX3 U634 ( .A(n1972), .Y(n1967) );
  CLKBUFX3 U635 ( .A(n1972), .Y(n1968) );
  CLKBUFX3 U636 ( .A(n1973), .Y(n1969) );
  CLKBUFX3 U637 ( .A(n1973), .Y(n1970) );
  CLKBUFX3 U638 ( .A(n1466), .Y(n1460) );
  CLKBUFX3 U639 ( .A(n1963), .Y(n1957) );
  CLKBUFX3 U640 ( .A(n1529), .Y(n1535) );
  CLKBUFX3 U641 ( .A(n1529), .Y(n1534) );
  CLKBUFX3 U642 ( .A(n2026), .Y(n2032) );
  CLKBUFX3 U643 ( .A(n2026), .Y(n2031) );
  CLKBUFX3 U644 ( .A(n1530), .Y(n1533) );
  CLKBUFX3 U645 ( .A(n1530), .Y(n1532) );
  CLKBUFX3 U646 ( .A(n1497), .Y(n1500) );
  CLKBUFX3 U647 ( .A(n1497), .Y(n1501) );
  CLKBUFX3 U648 ( .A(n1497), .Y(n1499) );
  CLKBUFX3 U649 ( .A(n1994), .Y(n1997) );
  CLKBUFX3 U650 ( .A(n2027), .Y(n2029) );
  CLKBUFX3 U651 ( .A(n1994), .Y(n1996) );
  CLKBUFX3 U652 ( .A(n2027), .Y(n2030) );
  CLKBUFX3 U653 ( .A(n1994), .Y(n1998) );
  CLKBUFX3 U654 ( .A(n1531), .Y(n1502) );
  CLKBUFX3 U655 ( .A(n1530), .Y(n1531) );
  CLKBUFX3 U656 ( .A(n2028), .Y(n1999) );
  CLKBUFX3 U657 ( .A(n2027), .Y(n2028) );
  CLKINVX1 U658 ( .A(n2253), .Y(n2364) );
  NAND2BX1 U659 ( .AN(n1951), .B(n1950), .Y(n1607) );
  MXI2X1 U660 ( .A(n1538), .B(n1539), .S0(n1952), .Y(ReadData2[1]) );
  MX4X1 U661 ( .A(n1615), .B(n1613), .C(n1614), .D(n1612), .S0(n1957), .S1(
        n1966), .Y(n1538) );
  MX4X1 U662 ( .A(n1611), .B(n1609), .C(n1610), .D(n1608), .S0(n1957), .S1(
        n1966), .Y(n1539) );
  NAND2BX1 U663 ( .AN(n1948), .B(n1947), .Y(n1615) );
  MXI2X1 U664 ( .A(n1540), .B(n1541), .S0(n1952), .Y(ReadData2[2]) );
  MX4X1 U665 ( .A(n1623), .B(n1621), .C(n1622), .D(n1620), .S0(n1958), .S1(
        n1966), .Y(n1540) );
  MX4X1 U666 ( .A(n1619), .B(n1617), .C(n1618), .D(n1616), .S0(n1958), .S1(
        n1966), .Y(n1541) );
  NAND2BX1 U667 ( .AN(n1945), .B(n1944), .Y(n1623) );
  MXI2X1 U668 ( .A(n1542), .B(n1543), .S0(n1952), .Y(ReadData2[3]) );
  MX4X1 U669 ( .A(n1631), .B(n1629), .C(n1630), .D(n1628), .S0(n1958), .S1(
        n1966), .Y(n1542) );
  MX4X1 U670 ( .A(n1627), .B(n1625), .C(n1626), .D(n1624), .S0(n1958), .S1(
        n1966), .Y(n1543) );
  NAND2BX1 U671 ( .AN(n1942), .B(n1941), .Y(n1631) );
  MXI2X1 U672 ( .A(n1544), .B(n1545), .S0(n1952), .Y(ReadData2[4]) );
  MX4X1 U673 ( .A(n1639), .B(n1637), .C(n1638), .D(n1636), .S0(n1958), .S1(
        n1966), .Y(n1544) );
  MX4X1 U674 ( .A(n1635), .B(n1633), .C(n1634), .D(n1632), .S0(n1958), .S1(
        n1966), .Y(n1545) );
  NAND2BX1 U675 ( .AN(n1939), .B(n1938), .Y(n1639) );
  MXI2X1 U676 ( .A(n1546), .B(n1547), .S0(n1952), .Y(ReadData2[5]) );
  MX4X1 U677 ( .A(n1647), .B(n1645), .C(n1646), .D(n1644), .S0(n1958), .S1(
        n1966), .Y(n1546) );
  MX4X1 U678 ( .A(n1643), .B(n1641), .C(n1642), .D(n1640), .S0(n1958), .S1(
        n1966), .Y(n1547) );
  NAND2BX1 U679 ( .AN(n1936), .B(n1935), .Y(n1647) );
  MXI2X1 U680 ( .A(n1548), .B(n1549), .S0(n1952), .Y(ReadData2[6]) );
  MX4X1 U681 ( .A(n1655), .B(n1653), .C(n1654), .D(n1652), .S0(n1958), .S1(
        n1967), .Y(n1548) );
  MX4X1 U682 ( .A(n1651), .B(n1649), .C(n1650), .D(n1648), .S0(n1958), .S1(
        n1967), .Y(n1549) );
  NAND2BX1 U683 ( .AN(n1933), .B(n1932), .Y(n1655) );
  MXI2X1 U684 ( .A(n1550), .B(n1551), .S0(n1952), .Y(ReadData2[7]) );
  MX4X1 U685 ( .A(n1663), .B(n1661), .C(n1662), .D(n1660), .S0(n1958), .S1(
        n1967), .Y(n1550) );
  MX4X1 U686 ( .A(n1659), .B(n1657), .C(n1658), .D(n1656), .S0(n1958), .S1(
        n1967), .Y(n1551) );
  NAND2BX1 U687 ( .AN(n1930), .B(n1929), .Y(n1663) );
  MXI2X1 U688 ( .A(n1552), .B(n1553), .S0(n1953), .Y(ReadData2[8]) );
  MX4X1 U689 ( .A(n1671), .B(n1669), .C(n1670), .D(n1668), .S0(n1959), .S1(
        n1967), .Y(n1552) );
  MX4X1 U690 ( .A(n1667), .B(n1665), .C(n1666), .D(n1664), .S0(n1959), .S1(
        n1967), .Y(n1553) );
  NAND2BX1 U691 ( .AN(n1927), .B(n1926), .Y(n1671) );
  MXI2X1 U692 ( .A(n1554), .B(n1555), .S0(n1953), .Y(ReadData2[9]) );
  MX4X1 U693 ( .A(n1679), .B(n1677), .C(n1678), .D(n1676), .S0(n1959), .S1(
        n1967), .Y(n1554) );
  MX4X1 U694 ( .A(n1675), .B(n1673), .C(n1674), .D(n1672), .S0(n1959), .S1(
        n1967), .Y(n1555) );
  NAND2BX1 U695 ( .AN(n1924), .B(n1923), .Y(n1679) );
  MXI2X1 U696 ( .A(n1556), .B(n1557), .S0(n1953), .Y(ReadData2[10]) );
  MX4X1 U697 ( .A(n1687), .B(n1685), .C(n1686), .D(n1684), .S0(n1959), .S1(
        n1967), .Y(n1556) );
  MX4X1 U698 ( .A(n1683), .B(n1681), .C(n1682), .D(n1680), .S0(n1959), .S1(
        n1967), .Y(n1557) );
  NAND2BX1 U699 ( .AN(n1921), .B(n1920), .Y(n1687) );
  MXI2X1 U700 ( .A(n1558), .B(n1559), .S0(n1953), .Y(ReadData2[11]) );
  MX4X1 U701 ( .A(n1695), .B(n1693), .C(n1694), .D(n1692), .S0(n1959), .S1(
        n1967), .Y(n1558) );
  MX4X1 U702 ( .A(n1691), .B(n1689), .C(n1690), .D(n1688), .S0(n1959), .S1(
        n1967), .Y(n1559) );
  NAND2BX1 U703 ( .AN(n1918), .B(n1917), .Y(n1695) );
  MXI2X1 U704 ( .A(n1560), .B(n1561), .S0(n1953), .Y(ReadData2[12]) );
  MX4X1 U705 ( .A(n1703), .B(n1701), .C(n1702), .D(n1700), .S0(n1959), .S1(
        n1968), .Y(n1560) );
  MX4X1 U706 ( .A(n1699), .B(n1697), .C(n1698), .D(n1696), .S0(n1959), .S1(
        n1967), .Y(n1561) );
  NAND2BX1 U707 ( .AN(n1915), .B(n1914), .Y(n1703) );
  MXI2X1 U708 ( .A(n1562), .B(n1563), .S0(n1953), .Y(ReadData2[13]) );
  MX4X1 U709 ( .A(n1711), .B(n1709), .C(n1710), .D(n1708), .S0(n1959), .S1(
        n1968), .Y(n1562) );
  MX4X1 U710 ( .A(n1707), .B(n1705), .C(n1706), .D(n1704), .S0(n1959), .S1(
        n1968), .Y(n1563) );
  NAND2BX1 U711 ( .AN(n1912), .B(n1911), .Y(n1711) );
  CLKINVX1 U712 ( .A(WriteData[28]), .Y(n2400) );
  CLKINVX1 U713 ( .A(WriteData[29]), .Y(n2399) );
  CLKINVX1 U714 ( .A(WriteData[30]), .Y(n2398) );
  CLKINVX1 U715 ( .A(WriteData[31]), .Y(n2397) );
  CLKINVX1 U716 ( .A(WriteData[0]), .Y(n2432) );
  CLKINVX1 U717 ( .A(WriteData[1]), .Y(n2427) );
  CLKINVX1 U718 ( .A(WriteData[2]), .Y(n2426) );
  CLKINVX1 U719 ( .A(WriteData[3]), .Y(n2425) );
  CLKINVX1 U720 ( .A(WriteData[4]), .Y(n2424) );
  CLKINVX1 U721 ( .A(WriteData[5]), .Y(n2423) );
  CLKINVX1 U722 ( .A(WriteData[6]), .Y(n2422) );
  CLKINVX1 U723 ( .A(WriteData[7]), .Y(n2421) );
  CLKINVX1 U724 ( .A(WriteData[8]), .Y(n2420) );
  CLKINVX1 U725 ( .A(WriteData[9]), .Y(n2419) );
  CLKINVX1 U726 ( .A(WriteData[10]), .Y(n2418) );
  CLKINVX1 U727 ( .A(WriteData[11]), .Y(n2417) );
  CLKINVX1 U728 ( .A(WriteData[12]), .Y(n2416) );
  CLKINVX1 U729 ( .A(WriteData[13]), .Y(n2415) );
  CLKINVX1 U730 ( .A(WriteData[14]), .Y(n2414) );
  CLKINVX1 U731 ( .A(WriteData[15]), .Y(n2413) );
  CLKINVX1 U732 ( .A(WriteData[16]), .Y(n2412) );
  CLKINVX1 U733 ( .A(WriteData[17]), .Y(n2411) );
  CLKINVX1 U734 ( .A(WriteData[18]), .Y(n2410) );
  CLKINVX1 U735 ( .A(WriteData[19]), .Y(n2409) );
  CLKINVX1 U736 ( .A(WriteData[20]), .Y(n2408) );
  CLKINVX1 U737 ( .A(WriteData[21]), .Y(n2407) );
  CLKINVX1 U738 ( .A(WriteData[22]), .Y(n2406) );
  CLKINVX1 U739 ( .A(WriteData[23]), .Y(n2405) );
  CLKINVX1 U740 ( .A(WriteData[24]), .Y(n2404) );
  CLKINVX1 U741 ( .A(WriteData[25]), .Y(n2403) );
  CLKINVX1 U742 ( .A(WriteData[26]), .Y(n2402) );
  CLKINVX1 U743 ( .A(WriteData[27]), .Y(n2401) );
  AND3X2 U744 ( .A(n53), .B(n2431), .C(WriteReg[4]), .Y(n65) );
  AND3X2 U745 ( .A(WriteReg[3]), .B(n53), .C(WriteReg[4]), .Y(n74) );
  CLKBUFX3 U746 ( .A(n1459), .Y(n1456) );
  CLKBUFX3 U747 ( .A(n1459), .Y(n1457) );
  CLKBUFX3 U748 ( .A(n1956), .Y(n1953) );
  CLKBUFX3 U749 ( .A(n1956), .Y(n1954) );
  CLKBUFX3 U750 ( .A(n1475), .Y(n1470) );
  CLKBUFX3 U751 ( .A(n1475), .Y(n1471) );
  CLKBUFX3 U752 ( .A(n1476), .Y(n1472) );
  CLKBUFX3 U753 ( .A(n1476), .Y(n1473) );
  CLKBUFX3 U754 ( .A(n1971), .Y(n1966) );
  CLKBUFX3 U755 ( .A(N20), .Y(n1971) );
  CLKBUFX3 U756 ( .A(rst_n), .Y(n2253) );
  CLKINVX1 U757 ( .A(WriteReg[3]), .Y(n2431) );
  CLKBUFX3 U758 ( .A(N19), .Y(n1994) );
  CLKBUFX3 U759 ( .A(N14), .Y(n1497) );
  CLKBUFX3 U760 ( .A(N16), .Y(n1466) );
  CLKBUFX3 U761 ( .A(N16), .Y(n1467) );
  CLKBUFX3 U762 ( .A(N16), .Y(n1468) );
  CLKBUFX3 U763 ( .A(N21), .Y(n1963) );
  CLKBUFX3 U764 ( .A(N20), .Y(n1972) );
  CLKBUFX3 U765 ( .A(N21), .Y(n1964) );
  CLKBUFX3 U766 ( .A(N21), .Y(n1965) );
  CLKBUFX3 U767 ( .A(N20), .Y(n1973) );
  CLKBUFX3 U768 ( .A(N13), .Y(n1530) );
  CLKBUFX3 U769 ( .A(N18), .Y(n2027) );
  CLKBUFX3 U770 ( .A(N13), .Y(n1529) );
  CLKBUFX3 U771 ( .A(N18), .Y(n2026) );
  MX4X1 U772 ( .A(n1106), .B(n1104), .C(n1105), .D(n1103), .S0(n1460), .S1(
        n1469), .Y(n4) );
  MX4X1 U773 ( .A(n1110), .B(n1108), .C(n1109), .D(n1107), .S0(n1460), .S1(
        n1469), .Y(n3) );
  MX4X1 U774 ( .A(n1114), .B(n1112), .C(n1113), .D(n1111), .S0(n1460), .S1(
        n1469), .Y(n6) );
  MX4X1 U775 ( .A(n1118), .B(n1116), .C(n1117), .D(n1115), .S0(n1460), .S1(
        n1469), .Y(n5) );
  MX4X1 U776 ( .A(n1162), .B(n1160), .C(n1161), .D(n1159), .S0(n1461), .S1(
        n1470), .Y(n18) );
  MX4X1 U777 ( .A(n1166), .B(n1164), .C(n1165), .D(n1163), .S0(n1461), .S1(
        n1470), .Y(n17) );
  MXI2X1 U778 ( .A(n19), .B(n20), .S0(n1456), .Y(ReadData1[8]) );
  MX4X1 U779 ( .A(n1170), .B(n1168), .C(n1169), .D(n1167), .S0(n1462), .S1(
        n1470), .Y(n20) );
  MX4X1 U780 ( .A(n1174), .B(n1172), .C(n1173), .D(n1171), .S0(n1462), .S1(
        n1470), .Y(n19) );
  MXI2X1 U781 ( .A(n9), .B(n10), .S0(n1455), .Y(ReadData1[3]) );
  MX4X1 U782 ( .A(n1130), .B(n1128), .C(n1129), .D(n1127), .S0(n1461), .S1(
        n1469), .Y(n10) );
  MX4X1 U783 ( .A(n1134), .B(n1132), .C(n1133), .D(n1131), .S0(n1461), .S1(
        n1469), .Y(n9) );
  MXI2X1 U784 ( .A(n7), .B(n8), .S0(n1455), .Y(ReadData1[2]) );
  MX4X1 U785 ( .A(n1122), .B(n1120), .C(n1121), .D(n1119), .S0(n1461), .S1(
        n1469), .Y(n8) );
  MX4X1 U786 ( .A(n1126), .B(n1124), .C(n1125), .D(n1123), .S0(n1461), .S1(
        n1469), .Y(n7) );
  NAND2BX1 U787 ( .AN(n1448), .B(n1447), .Y(n1126) );
  OAI22XL U788 ( .A0(n1496), .A1(n1524), .B0(n1492), .B1(\register[1][2] ), 
        .Y(n1448) );
  NAND2BX1 U789 ( .AN(n1433), .B(n1432), .Y(n1166) );
  MXI2X1 U790 ( .A(n2372), .B(n1431), .S0(n1527), .Y(n1432) );
  OAI22XL U791 ( .A0(n1495), .A1(n1524), .B0(n1492), .B1(\register[1][7] ), 
        .Y(n1433) );
  NAND2BX1 U792 ( .AN(n1454), .B(n1453), .Y(n1110) );
  MXI2X1 U793 ( .A(n2365), .B(n1452), .S0(n1528), .Y(n1453) );
  OAI22XL U794 ( .A0(n1496), .A1(n1525), .B0(n1491), .B1(\register[1][0] ), 
        .Y(n1454) );
  OAI22XL U795 ( .A0(n1993), .A1(n2021), .B0(n1989), .B1(\register[1][2] ), 
        .Y(n1945) );
  OAI22XL U796 ( .A0(n1993), .A1(n2021), .B0(n1989), .B1(\register[1][3] ), 
        .Y(n1942) );
  OAI22XL U797 ( .A0(n1993), .A1(n2021), .B0(n1989), .B1(\register[1][4] ), 
        .Y(n1939) );
  OAI22XL U798 ( .A0(n1992), .A1(n2021), .B0(n1989), .B1(\register[1][5] ), 
        .Y(n1936) );
  OAI22XL U799 ( .A0(n1993), .A1(n2021), .B0(n1989), .B1(\register[1][6] ), 
        .Y(n1933) );
  OAI22XL U800 ( .A0(n1992), .A1(n2021), .B0(n1989), .B1(\register[1][7] ), 
        .Y(n1930) );
  OAI22XL U801 ( .A0(n1992), .A1(n2021), .B0(n1989), .B1(\register[1][8] ), 
        .Y(n1927) );
  MXI2X1 U802 ( .A(n2365), .B(n1949), .S0(n2025), .Y(n1950) );
  NOR2BX1 U803 ( .AN(n1987), .B(\register[3][0] ), .Y(n1949) );
  MXI2X1 U804 ( .A(n2366), .B(n1946), .S0(n2025), .Y(n1947) );
  NOR2BX1 U805 ( .AN(n1988), .B(\register[3][1] ), .Y(n1946) );
  MXI2X1 U806 ( .A(n2367), .B(n1943), .S0(n2025), .Y(n1944) );
  NOR2BX1 U807 ( .AN(n1988), .B(\register[3][2] ), .Y(n1943) );
  MXI2X1 U808 ( .A(n2368), .B(n1940), .S0(n2025), .Y(n1941) );
  NOR2BX1 U809 ( .AN(n1988), .B(\register[3][3] ), .Y(n1940) );
  MXI2X1 U810 ( .A(n2369), .B(n1937), .S0(n2025), .Y(n1938) );
  NOR2BX1 U811 ( .AN(n1988), .B(\register[3][4] ), .Y(n1937) );
  MXI2X1 U812 ( .A(n2370), .B(n1934), .S0(n2025), .Y(n1935) );
  NOR2BX1 U813 ( .AN(n1988), .B(\register[3][5] ), .Y(n1934) );
  MXI2X1 U814 ( .A(n2371), .B(n1931), .S0(n2025), .Y(n1932) );
  NOR2BX1 U815 ( .AN(n1988), .B(\register[3][6] ), .Y(n1931) );
  MXI2X1 U816 ( .A(n2372), .B(n1928), .S0(n2024), .Y(n1929) );
  NOR2BX1 U817 ( .AN(n1988), .B(\register[3][7] ), .Y(n1928) );
  MXI2X1 U818 ( .A(n2373), .B(n1925), .S0(n2025), .Y(n1926) );
  NOR2BX1 U819 ( .AN(n1988), .B(\register[3][8] ), .Y(n1925) );
  MX4X1 U820 ( .A(n1138), .B(n1136), .C(n1137), .D(n1135), .S0(n1461), .S1(
        n1469), .Y(n12) );
  MX4X1 U821 ( .A(n1142), .B(n1140), .C(n1141), .D(n1139), .S0(n1461), .S1(
        n1469), .Y(n11) );
  MX4X1 U822 ( .A(n1146), .B(n1144), .C(n1145), .D(n1143), .S0(n1461), .S1(
        n1469), .Y(n14) );
  MX4X1 U823 ( .A(n1150), .B(n1148), .C(n1149), .D(n1147), .S0(n1461), .S1(
        n1469), .Y(n13) );
  MX4X1 U824 ( .A(n1154), .B(n1152), .C(n1153), .D(n1151), .S0(n1461), .S1(
        n1470), .Y(n16) );
  MX4X1 U825 ( .A(n1158), .B(n1156), .C(n1157), .D(n1155), .S0(n1461), .S1(
        n1470), .Y(n15) );
  NAND2BX1 U826 ( .AN(n1445), .B(n1444), .Y(n1134) );
  OAI22XL U827 ( .A0(n1496), .A1(n1524), .B0(n1492), .B1(\register[1][3] ), 
        .Y(n1445) );
  NAND2BX1 U828 ( .AN(n1442), .B(n1441), .Y(n1142) );
  MXI2X1 U829 ( .A(n2369), .B(n1440), .S0(n1528), .Y(n1441) );
  OAI22XL U830 ( .A0(n1496), .A1(n1524), .B0(n1492), .B1(\register[1][4] ), 
        .Y(n1442) );
  NAND2BX1 U831 ( .AN(n1439), .B(n1438), .Y(n1150) );
  MXI2X1 U832 ( .A(n2370), .B(n1437), .S0(n1528), .Y(n1438) );
  OAI22XL U833 ( .A0(n1495), .A1(n1524), .B0(n1492), .B1(\register[1][5] ), 
        .Y(n1439) );
  NAND2BX1 U834 ( .AN(n1436), .B(n1435), .Y(n1158) );
  MXI2X1 U835 ( .A(n2371), .B(n1434), .S0(n1528), .Y(n1435) );
  OAI22XL U836 ( .A0(n1496), .A1(n1524), .B0(n1492), .B1(\register[1][6] ), 
        .Y(n1436) );
  NAND2BX1 U837 ( .AN(n1430), .B(n1429), .Y(n1174) );
  OAI22XL U838 ( .A0(n1495), .A1(n1524), .B0(n1492), .B1(\register[1][8] ), 
        .Y(n1430) );
  NAND2BX1 U839 ( .AN(n1451), .B(n1450), .Y(n1118) );
  MXI2X1 U840 ( .A(n2366), .B(n1449), .S0(n1528), .Y(n1450) );
  OAI22XL U841 ( .A0(n1496), .A1(n1524), .B0(n1492), .B1(\register[1][1] ), 
        .Y(n1451) );
  MXI4X1 U842 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n2014), .S1(n1984), .Y(
        n1602) );
  MXI4X1 U843 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n2014), .S1(n1985), .Y(
        n1606) );
  MXI4X1 U844 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n2015), .S1(n1985), .Y(
        n1610) );
  MXI4X1 U845 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n2015), .S1(n1985), .Y(
        n1614) );
  MXI4X1 U846 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n2015), .S1(n1985), .Y(
        n1618) );
  MXI4X1 U847 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n2015), .S1(n1985), .Y(
        n1622) );
  MXI4X1 U848 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n2015), .S1(n1985), .Y(
        n1626) );
  MXI4X1 U849 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n2016), .S1(n1985), .Y(
        n1630) );
  MXI4X1 U850 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n2016), .S1(n1985), .Y(
        n1634) );
  MXI4X1 U851 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n2016), .S1(n1985), .Y(
        n1638) );
  MXI4X1 U852 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n2016), .S1(n1985), .Y(
        n1642) );
  MXI4X1 U853 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n2016), .S1(n1986), .Y(
        n1646) );
  MXI4X1 U854 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n2017), .S1(n1986), .Y(
        n1650) );
  MXI4X1 U855 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n2017), .S1(n1986), .Y(
        n1654) );
  MXI4X1 U856 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n2017), .S1(n1986), .Y(
        n1658) );
  MXI4X1 U857 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n2017), .S1(n1986), .Y(
        n1662) );
  MXI4X1 U858 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n2018), .S1(n1987), .Y(
        n1666) );
  MXI4X1 U859 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n2018), .S1(n1987), .Y(
        n1670) );
  MXI4X1 U860 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n2014), .S1(n1985), .Y(
        n1603) );
  MXI4X1 U861 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n2015), .S1(n1985), .Y(
        n1611) );
  MXI4X1 U862 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n2015), .S1(n1985), .Y(
        n1619) );
  MXI4X1 U863 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n2015), .S1(n1985), .Y(
        n1627) );
  MXI4X1 U864 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n2016), .S1(n1985), .Y(
        n1635) );
  MXI4X1 U865 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n2016), .S1(n1985), .Y(
        n1643) );
  MXI4X1 U866 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n2017), .S1(n1986), .Y(
        n1651) );
  MXI4X1 U867 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n2017), .S1(n1986), .Y(
        n1659) );
  MXI4X1 U868 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n2018), .S1(n1987), .Y(
        n1667) );
  MXI4X1 U869 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n2014), .S1(n1984), .Y(
        n1600) );
  MXI4X1 U870 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n2014), .S1(n1985), .Y(
        n1604) );
  MXI4X1 U871 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n2014), .S1(n1985), .Y(
        n1608) );
  MXI4X1 U872 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n2015), .S1(n1985), .Y(
        n1612) );
  MXI4X1 U873 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n2015), .S1(n1985), .Y(
        n1616) );
  MXI4X1 U874 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n2015), .S1(n1985), .Y(
        n1620) );
  MXI4X1 U875 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n2015), .S1(n1985), .Y(
        n1624) );
  MXI4X1 U876 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n2016), .S1(n1985), .Y(
        n1628) );
  MXI4X1 U877 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n2016), .S1(n1985), .Y(
        n1632) );
  MXI4X1 U878 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n2016), .S1(n1985), .Y(
        n1636) );
  MXI4X1 U879 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n2016), .S1(n1985), .Y(
        n1640) );
  MXI4X1 U880 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n2016), .S1(n1985), .Y(
        n1644) );
  MXI4X1 U881 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n2017), .S1(n1986), .Y(
        n1648) );
  MXI4X1 U882 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n2017), .S1(n1986), .Y(
        n1652) );
  MXI4X1 U883 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n2017), .S1(n1986), .Y(
        n1656) );
  MXI4X1 U884 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n2017), .S1(n1986), .Y(
        n1660) );
  MXI4X1 U885 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n2017), .S1(n1987), .Y(
        n1664) );
  MXI4X1 U886 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n2018), .S1(n1987), .Y(
        n1668) );
  MXI4X1 U887 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n2014), .S1(n1984), .Y(
        n1601) );
  MXI4X1 U888 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n2014), .S1(n1985), .Y(
        n1605) );
  MXI4X1 U889 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n2015), .S1(n1985), .Y(
        n1609) );
  MXI4X1 U890 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n2015), .S1(n1985), .Y(
        n1613) );
  MXI4X1 U891 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n2015), .S1(n1985), .Y(
        n1617) );
  MXI4X1 U892 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n2015), .S1(n1985), .Y(
        n1621) );
  MXI4X1 U893 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n2015), .S1(n1985), .Y(
        n1625) );
  MXI4X1 U894 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n2016), .S1(n1985), .Y(
        n1629) );
  MXI4X1 U895 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n2016), .S1(n1985), .Y(
        n1633) );
  MXI4X1 U896 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n2016), .S1(n1985), .Y(
        n1637) );
  MXI4X1 U897 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n2016), .S1(n1985), .Y(
        n1641) );
  MXI4X1 U898 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n2016), .S1(n1986), .Y(
        n1645) );
  MXI4X1 U899 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n2017), .S1(n1986), .Y(
        n1649) );
  MXI4X1 U900 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n2017), .S1(n1986), .Y(
        n1653) );
  MXI4X1 U901 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n2017), .S1(n1986), .Y(
        n1657) );
  MXI4X1 U902 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n2017), .S1(n1986), .Y(
        n1661) );
  MXI4X1 U903 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n2017), .S1(n1987), .Y(
        n1665) );
  MXI4X1 U904 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n2018), .S1(n1987), .Y(
        n1669) );
  MX4X1 U905 ( .A(n1218), .B(n1216), .C(n1217), .D(n1215), .S0(n1463), .S1(
        n1471), .Y(n32) );
  MX4X1 U906 ( .A(n1222), .B(n1220), .C(n1221), .D(n1219), .S0(n1463), .S1(
        n1471), .Y(n31) );
  MX4X1 U907 ( .A(n1234), .B(n1232), .C(n1233), .D(n1231), .S0(n1463), .S1(
        n1471), .Y(n36) );
  MX4X1 U908 ( .A(n1238), .B(n1236), .C(n1237), .D(n1235), .S0(n1463), .S1(
        n1471), .Y(n35) );
  MX4X1 U909 ( .A(n1242), .B(n1240), .C(n1241), .D(n1239), .S0(n1463), .S1(
        n1471), .Y(n1074) );
  MX4X1 U910 ( .A(n1246), .B(n1244), .C(n1245), .D(n1243), .S0(n1463), .S1(
        n1471), .Y(n37) );
  MXI4X1 U911 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1239) );
  MX4X1 U912 ( .A(n1282), .B(n1280), .C(n1281), .D(n1279), .S0(n1464), .S1(
        n1472), .Y(n1084) );
  MX4X1 U913 ( .A(n1286), .B(n1284), .C(n1285), .D(n1283), .S0(n1464), .S1(
        n1472), .Y(n1083) );
  MXI4X1 U914 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1279) );
  MXI2X1 U915 ( .A(n1075), .B(n1076), .S0(n1456), .Y(ReadData1[18]) );
  MX4X1 U916 ( .A(n1250), .B(n1248), .C(n1249), .D(n1247), .S0(n1463), .S1(
        n1471), .Y(n1076) );
  MX4X1 U917 ( .A(n1254), .B(n1252), .C(n1253), .D(n1251), .S0(n1463), .S1(
        n1471), .Y(n1075) );
  MXI4X1 U918 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1511), .S1(n1485), 
        .Y(n1247) );
  MXI2X1 U919 ( .A(n21), .B(n22), .S0(n1456), .Y(ReadData1[9]) );
  MX4X1 U920 ( .A(n1178), .B(n1176), .C(n1177), .D(n1175), .S0(n1462), .S1(
        n1470), .Y(n22) );
  MX4X1 U921 ( .A(n1182), .B(n1180), .C(n1181), .D(n1179), .S0(n1462), .S1(
        n1470), .Y(n21) );
  MXI2X1 U922 ( .A(n1077), .B(n1078), .S0(n1456), .Y(ReadData1[19]) );
  MX4X1 U923 ( .A(n1258), .B(n1256), .C(n1257), .D(n1255), .S0(n1463), .S1(
        n1472), .Y(n1078) );
  MX4X1 U924 ( .A(n1262), .B(n1260), .C(n1261), .D(n1259), .S0(n1463), .S1(
        n1472), .Y(n1077) );
  MXI4X1 U925 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1255) );
  MXI2X1 U926 ( .A(n25), .B(n26), .S0(n1456), .Y(ReadData1[11]) );
  MX4X1 U927 ( .A(n1194), .B(n1192), .C(n1193), .D(n1191), .S0(n1462), .S1(
        n1470), .Y(n26) );
  MX4X1 U928 ( .A(n1198), .B(n1196), .C(n1197), .D(n1195), .S0(n1462), .S1(
        n1470), .Y(n25) );
  MXI2X1 U929 ( .A(n29), .B(n30), .S0(n1456), .Y(ReadData1[13]) );
  MX4X1 U930 ( .A(n1210), .B(n1208), .C(n1209), .D(n1207), .S0(n1462), .S1(
        n1471), .Y(n30) );
  MX4X1 U931 ( .A(n1214), .B(n1212), .C(n1213), .D(n1211), .S0(n1462), .S1(
        n1471), .Y(n29) );
  MXI2X1 U932 ( .A(n1081), .B(n1082), .S0(n1457), .Y(ReadData1[21]) );
  MX4X1 U933 ( .A(n1274), .B(n1272), .C(n1273), .D(n1271), .S0(n1464), .S1(
        n1472), .Y(n1082) );
  MX4X1 U934 ( .A(n1278), .B(n1276), .C(n1277), .D(n1275), .S0(n1464), .S1(
        n1472), .Y(n1081) );
  MXI4X1 U935 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1513), .S1(n1485), 
        .Y(n1271) );
  MXI2X1 U936 ( .A(n23), .B(n24), .S0(n1456), .Y(ReadData1[10]) );
  MX4X1 U937 ( .A(n1186), .B(n1184), .C(n1185), .D(n1183), .S0(n1462), .S1(
        n1470), .Y(n24) );
  MX4X1 U938 ( .A(n1190), .B(n1188), .C(n1189), .D(n1187), .S0(n1462), .S1(
        n1470), .Y(n23) );
  MXI2X1 U939 ( .A(n27), .B(n28), .S0(n1456), .Y(ReadData1[12]) );
  MX4X1 U940 ( .A(n1202), .B(n1200), .C(n1201), .D(n1199), .S0(n1462), .S1(
        n1470), .Y(n28) );
  MX4X1 U941 ( .A(n1206), .B(n1204), .C(n1205), .D(n1203), .S0(n1462), .S1(
        n1471), .Y(n27) );
  MXI2X1 U942 ( .A(n1079), .B(n1080), .S0(n1457), .Y(ReadData1[20]) );
  MX4X1 U943 ( .A(n1266), .B(n1264), .C(n1265), .D(n1263), .S0(n1464), .S1(
        n1472), .Y(n1080) );
  MX4X1 U944 ( .A(n1270), .B(n1268), .C(n1269), .D(n1267), .S0(n1464), .S1(
        n1472), .Y(n1079) );
  MXI4X1 U945 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1263) );
  MXI2X1 U946 ( .A(n33), .B(n34), .S0(n1456), .Y(ReadData1[15]) );
  MX4X1 U947 ( .A(n1226), .B(n1224), .C(n1225), .D(n1223), .S0(n1463), .S1(
        n1471), .Y(n34) );
  MX4X1 U948 ( .A(n1230), .B(n1228), .C(n1229), .D(n1227), .S0(n1463), .S1(
        n1471), .Y(n33) );
  MXI4X1 U949 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1523), .S1(n1489), 
        .Y(n1223) );
  OAI22XL U950 ( .A0(n1992), .A1(n2021), .B0(n1989), .B1(\register[1][9] ), 
        .Y(n1924) );
  OAI22XL U951 ( .A0(n1992), .A1(n2021), .B0(n1989), .B1(\register[1][10] ), 
        .Y(n1921) );
  OAI22XL U952 ( .A0(n1991), .A1(n2021), .B0(n1989), .B1(\register[1][11] ), 
        .Y(n1918) );
  OAI22XL U953 ( .A0(n1991), .A1(n2021), .B0(n1990), .B1(\register[1][12] ), 
        .Y(n1915) );
  OAI22XL U954 ( .A0(n1991), .A1(n2022), .B0(n1989), .B1(\register[1][13] ), 
        .Y(n1912) );
  MXI2X1 U955 ( .A(n2374), .B(n1922), .S0(n2024), .Y(n1923) );
  NOR2BX1 U956 ( .AN(n1988), .B(\register[3][9] ), .Y(n1922) );
  MXI2X1 U957 ( .A(n2375), .B(n1919), .S0(n2024), .Y(n1920) );
  NOR2BX1 U958 ( .AN(n1988), .B(\register[3][10] ), .Y(n1919) );
  MXI2X1 U959 ( .A(n2376), .B(n1916), .S0(n2024), .Y(n1917) );
  NOR2BX1 U960 ( .AN(n1988), .B(\register[3][11] ), .Y(n1916) );
  MXI2X1 U961 ( .A(n2377), .B(n1913), .S0(n2024), .Y(n1914) );
  NOR2BX1 U962 ( .AN(n1988), .B(\register[3][12] ), .Y(n1913) );
  MXI2X1 U963 ( .A(n2378), .B(n1910), .S0(n2024), .Y(n1911) );
  NOR2BX1 U964 ( .AN(n1988), .B(\register[3][13] ), .Y(n1910) );
  MXI2X1 U965 ( .A(n1564), .B(n1565), .S0(n1953), .Y(ReadData2[14]) );
  MX4X1 U966 ( .A(n1715), .B(n1713), .C(n1714), .D(n1712), .S0(n1960), .S1(
        n1968), .Y(n1565) );
  MX4X1 U967 ( .A(n1719), .B(n1717), .C(n1718), .D(n1716), .S0(n1960), .S1(
        n1968), .Y(n1564) );
  MXI4X1 U968 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1712) );
  MXI2X1 U969 ( .A(n1566), .B(n1567), .S0(n1953), .Y(ReadData2[15]) );
  MX4X1 U970 ( .A(n1723), .B(n1721), .C(n1722), .D(n1720), .S0(n1960), .S1(
        n1968), .Y(n1567) );
  MX4X1 U971 ( .A(n1727), .B(n1725), .C(n1726), .D(n1724), .S0(n1960), .S1(
        n1968), .Y(n1566) );
  MXI4X1 U972 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n2020), .S1(n1986), 
        .Y(n1720) );
  MXI2X1 U973 ( .A(n1568), .B(n1569), .S0(n1953), .Y(ReadData2[16]) );
  MX4X1 U974 ( .A(n1731), .B(n1729), .C(n1730), .D(n1728), .S0(n1960), .S1(
        n1968), .Y(n1569) );
  MX4X1 U975 ( .A(n1735), .B(n1733), .C(n1734), .D(n1732), .S0(n1960), .S1(
        n1968), .Y(n1568) );
  MXI4X1 U976 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n2008), .S1(n1981), 
        .Y(n1728) );
  MXI2X1 U977 ( .A(n1570), .B(n1571), .S0(n1953), .Y(ReadData2[17]) );
  MX4X1 U978 ( .A(n1739), .B(n1737), .C(n1738), .D(n1736), .S0(n1960), .S1(
        n1968), .Y(n1571) );
  MX4X1 U979 ( .A(n1743), .B(n1741), .C(n1742), .D(n1740), .S0(n1960), .S1(
        n1968), .Y(n1570) );
  MXI4X1 U980 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1736) );
  MXI2X1 U981 ( .A(n1572), .B(n1573), .S0(n1953), .Y(ReadData2[18]) );
  MX4X1 U982 ( .A(n1747), .B(n1745), .C(n1746), .D(n1744), .S0(n1960), .S1(
        n1968), .Y(n1573) );
  MX4X1 U983 ( .A(n1751), .B(n1749), .C(n1750), .D(n1748), .S0(n1960), .S1(
        n1968), .Y(n1572) );
  MXI4X1 U984 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n2008), .S1(n1982), 
        .Y(n1744) );
  MXI2X1 U985 ( .A(n1574), .B(n1575), .S0(n1953), .Y(ReadData2[19]) );
  MX4X1 U986 ( .A(n1755), .B(n1753), .C(n1754), .D(n1752), .S0(n1960), .S1(
        n1969), .Y(n1575) );
  MX4X1 U987 ( .A(n1759), .B(n1757), .C(n1758), .D(n1756), .S0(n1960), .S1(
        n1969), .Y(n1574) );
  MXI4X1 U988 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1752) );
  MXI2X1 U989 ( .A(n1576), .B(n1577), .S0(n1954), .Y(ReadData2[20]) );
  MX4X1 U990 ( .A(n1763), .B(n1761), .C(n1762), .D(n1760), .S0(n1961), .S1(
        n1969), .Y(n1577) );
  MX4X1 U991 ( .A(n1767), .B(n1765), .C(n1766), .D(n1764), .S0(n1961), .S1(
        n1969), .Y(n1576) );
  MXI4X1 U992 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1760) );
  MXI2X1 U993 ( .A(n1578), .B(n1579), .S0(n1954), .Y(ReadData2[21]) );
  MX4X1 U994 ( .A(n1771), .B(n1769), .C(n1770), .D(n1768), .S0(n1961), .S1(
        n1969), .Y(n1579) );
  MX4X1 U995 ( .A(n1775), .B(n1773), .C(n1774), .D(n1772), .S0(n1961), .S1(
        n1969), .Y(n1578) );
  MXI4X1 U996 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n2010), .S1(n1982), 
        .Y(n1768) );
  MXI2X1 U997 ( .A(n1580), .B(n1581), .S0(n1954), .Y(ReadData2[22]) );
  MX4X1 U998 ( .A(n1779), .B(n1777), .C(n1778), .D(n1776), .S0(n1961), .S1(
        n1969), .Y(n1581) );
  MX4X1 U999 ( .A(n1783), .B(n1781), .C(n1782), .D(n1780), .S0(n1961), .S1(
        n1969), .Y(n1580) );
  MXI4X1 U1000 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1776) );
  MXI2X1 U1001 ( .A(n1582), .B(n1583), .S0(n1954), .Y(ReadData2[23]) );
  MX4X1 U1002 ( .A(n1787), .B(n1785), .C(n1786), .D(n1784), .S0(n1961), .S1(
        n1969), .Y(n1583) );
  MX4X1 U1003 ( .A(n1791), .B(n1789), .C(n1790), .D(n1788), .S0(n1961), .S1(
        n1969), .Y(n1582) );
  MXI4X1 U1004 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n2010), .S1(n1983), 
        .Y(n1784) );
  MXI2X1 U1005 ( .A(n1584), .B(n1585), .S0(n1954), .Y(ReadData2[24]) );
  MX4X1 U1006 ( .A(n1795), .B(n1793), .C(n1794), .D(n1792), .S0(n1961), .S1(
        n1969), .Y(n1585) );
  MX4X1 U1007 ( .A(n1799), .B(n1797), .C(n1798), .D(n1796), .S0(n1961), .S1(
        n1969), .Y(n1584) );
  MXI4X1 U1008 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1792) );
  MXI2X1 U1009 ( .A(n1586), .B(n1587), .S0(n1954), .Y(ReadData2[25]) );
  MX4X1 U1010 ( .A(n1803), .B(n1801), .C(n1802), .D(n1800), .S0(n1961), .S1(
        n1969), .Y(n1587) );
  MX4X1 U1011 ( .A(n1807), .B(n1805), .C(n1806), .D(n1804), .S0(n1961), .S1(
        n1970), .Y(n1586) );
  MXI4X1 U1012 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n2011), .S1(n1983), 
        .Y(n1800) );
  MXI2X1 U1013 ( .A(n1588), .B(n1589), .S0(n1954), .Y(ReadData2[26]) );
  MX4X1 U1014 ( .A(n1811), .B(n1809), .C(n1810), .D(n1808), .S0(n1962), .S1(
        n1970), .Y(n1589) );
  MX4X1 U1015 ( .A(n1815), .B(n1813), .C(n1814), .D(n1812), .S0(n1962), .S1(
        n1970), .Y(n1588) );
  MXI4X1 U1016 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1808) );
  MXI2X1 U1017 ( .A(n1590), .B(n1591), .S0(n1954), .Y(ReadData2[27]) );
  MX4X1 U1018 ( .A(n1819), .B(n1817), .C(n1818), .D(n1816), .S0(n1962), .S1(
        n1970), .Y(n1591) );
  MX4X1 U1019 ( .A(n1823), .B(n1821), .C(n1822), .D(n1820), .S0(n1962), .S1(
        n1970), .Y(n1590) );
  MXI4X1 U1020 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1816) );
  MXI2X1 U1021 ( .A(n1592), .B(n1593), .S0(n1954), .Y(ReadData2[28]) );
  MX4X1 U1022 ( .A(n1827), .B(n1825), .C(n1826), .D(n1824), .S0(n1962), .S1(
        n1970), .Y(n1593) );
  MX4X1 U1023 ( .A(n1831), .B(n1829), .C(n1830), .D(n1828), .S0(n1962), .S1(
        n1970), .Y(n1592) );
  MXI4X1 U1024 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1824) );
  MXI2X1 U1025 ( .A(n1594), .B(n1595), .S0(n1954), .Y(ReadData2[29]) );
  MX4X1 U1026 ( .A(n1835), .B(n1833), .C(n1834), .D(n1832), .S0(n1962), .S1(
        n1970), .Y(n1595) );
  MX4X1 U1027 ( .A(n1839), .B(n1837), .C(n1838), .D(n1836), .S0(n1962), .S1(
        n1970), .Y(n1594) );
  MXI4X1 U1028 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1832) );
  MXI2X1 U1029 ( .A(n1596), .B(n1597), .S0(n1954), .Y(ReadData2[30]) );
  MX4X1 U1030 ( .A(n1843), .B(n1841), .C(n1842), .D(n1840), .S0(n1962), .S1(
        n1970), .Y(n1597) );
  MX4X1 U1031 ( .A(n1847), .B(n1845), .C(n1846), .D(n1844), .S0(n1962), .S1(
        n1970), .Y(n1596) );
  MXI4X1 U1032 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n2013), .S1(n1984), 
        .Y(n1840) );
  MXI2X1 U1033 ( .A(n1598), .B(n1599), .S0(n1954), .Y(ReadData2[31]) );
  MX4X1 U1034 ( .A(n1851), .B(n1849), .C(n1850), .D(n1848), .S0(n1962), .S1(
        n1970), .Y(n1599) );
  MX4X1 U1035 ( .A(n1855), .B(n1853), .C(n1854), .D(n1852), .S0(n1962), .S1(
        n1970), .Y(n1598) );
  MXI4X1 U1036 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n2014), .S1(n1984), 
        .Y(n1848) );
  OAI2BB2XL U1037 ( .B0(n2128), .B1(n2245), .A0N(\register[2][0] ), .A1N(n2247), .Y(n114) );
  OAI2BB2XL U1038 ( .B0(n2125), .B1(n2245), .A0N(\register[2][1] ), .A1N(n2248), .Y(n115) );
  OAI2BB2XL U1039 ( .B0(n2122), .B1(n2245), .A0N(\register[2][2] ), .A1N(n2248), .Y(n116) );
  OAI2BB2XL U1040 ( .B0(n2119), .B1(n2245), .A0N(\register[2][3] ), .A1N(n2248), .Y(n117) );
  OAI2BB2XL U1041 ( .B0(n2116), .B1(n2245), .A0N(\register[2][4] ), .A1N(n2248), .Y(n118) );
  OAI2BB2XL U1042 ( .B0(n2113), .B1(n2245), .A0N(\register[2][5] ), .A1N(n2248), .Y(n119) );
  OAI2BB2XL U1043 ( .B0(n2110), .B1(n2245), .A0N(\register[2][6] ), .A1N(n2248), .Y(n120) );
  OAI2BB2XL U1044 ( .B0(n2107), .B1(n2245), .A0N(\register[2][7] ), .A1N(n2248), .Y(n121) );
  OAI2BB2XL U1045 ( .B0(n2104), .B1(n2246), .A0N(\register[2][8] ), .A1N(n2248), .Y(n122) );
  OAI2BB2XL U1046 ( .B0(n2101), .B1(n2246), .A0N(\register[2][9] ), .A1N(n2248), .Y(n123) );
  OAI2BB2XL U1047 ( .B0(n2098), .B1(n2246), .A0N(\register[2][10] ), .A1N(
        n2248), .Y(n124) );
  OAI2BB2XL U1048 ( .B0(n2095), .B1(n2246), .A0N(\register[2][11] ), .A1N(
        n2248), .Y(n125) );
  OAI2BB2XL U1049 ( .B0(n2092), .B1(n2246), .A0N(\register[2][12] ), .A1N(
        n2248), .Y(n126) );
  OAI2BB2XL U1050 ( .B0(n2089), .B1(n2246), .A0N(\register[2][13] ), .A1N(
        n2248), .Y(n127) );
  OAI2BB2XL U1051 ( .B0(n2086), .B1(n2246), .A0N(\register[2][14] ), .A1N(
        n2248), .Y(n128) );
  OAI2BB2XL U1052 ( .B0(n2083), .B1(n2246), .A0N(\register[2][15] ), .A1N(
        n2248), .Y(n129) );
  OAI2BB2XL U1053 ( .B0(n2080), .B1(n2247), .A0N(\register[2][16] ), .A1N(
        n2248), .Y(n130) );
  OAI2BB2XL U1054 ( .B0(n2077), .B1(n2247), .A0N(\register[2][17] ), .A1N(
        n2248), .Y(n131) );
  OAI2BB2XL U1055 ( .B0(n2074), .B1(n2246), .A0N(\register[2][18] ), .A1N(
        n2248), .Y(n132) );
  OAI2BB2XL U1056 ( .B0(n2071), .B1(n2247), .A0N(\register[2][19] ), .A1N(
        n2248), .Y(n133) );
  OAI2BB2XL U1057 ( .B0(n2068), .B1(n2247), .A0N(\register[2][20] ), .A1N(
        n2248), .Y(n134) );
  OAI2BB2XL U1058 ( .B0(n2065), .B1(n2247), .A0N(\register[2][21] ), .A1N(
        n2247), .Y(n135) );
  OAI2BB2XL U1059 ( .B0(n2062), .B1(n2247), .A0N(\register[2][22] ), .A1N(
        n2247), .Y(n136) );
  OAI2BB2XL U1060 ( .B0(n2059), .B1(n2247), .A0N(\register[2][23] ), .A1N(
        n2247), .Y(n137) );
  OAI2BB2XL U1061 ( .B0(n2056), .B1(n2247), .A0N(\register[2][24] ), .A1N(
        n2247), .Y(n138) );
  OAI2BB2XL U1062 ( .B0(n2053), .B1(n2246), .A0N(\register[2][25] ), .A1N(
        n2247), .Y(n139) );
  OAI2BB2XL U1063 ( .B0(n2050), .B1(n2246), .A0N(\register[2][26] ), .A1N(
        n2247), .Y(n140) );
  OAI2BB2XL U1064 ( .B0(n2047), .B1(n2246), .A0N(\register[2][27] ), .A1N(
        n2247), .Y(n141) );
  OAI2BB2XL U1065 ( .B0(n2044), .B1(n2245), .A0N(\register[2][28] ), .A1N(
        n2247), .Y(n142) );
  OAI2BB2XL U1066 ( .B0(n2041), .B1(n2245), .A0N(\register[2][29] ), .A1N(
        n2247), .Y(n143) );
  OAI2BB2XL U1067 ( .B0(n2038), .B1(n2245), .A0N(\register[2][30] ), .A1N(
        n2247), .Y(n144) );
  OAI2BB2XL U1068 ( .B0(n2035), .B1(n2245), .A0N(\register[2][31] ), .A1N(
        n2247), .Y(n145) );
  OAI2BB2XL U1069 ( .B0(n2128), .B1(n2241), .A0N(\register[3][0] ), .A1N(n2243), .Y(n146) );
  OAI2BB2XL U1070 ( .B0(n2125), .B1(n2241), .A0N(\register[3][1] ), .A1N(n2244), .Y(n147) );
  OAI2BB2XL U1071 ( .B0(n2122), .B1(n2241), .A0N(\register[3][2] ), .A1N(n2244), .Y(n148) );
  OAI2BB2XL U1072 ( .B0(n2119), .B1(n2241), .A0N(\register[3][3] ), .A1N(n2244), .Y(n149) );
  OAI2BB2XL U1073 ( .B0(n2116), .B1(n2241), .A0N(\register[3][4] ), .A1N(n2244), .Y(n150) );
  OAI2BB2XL U1074 ( .B0(n2113), .B1(n2241), .A0N(\register[3][5] ), .A1N(n2244), .Y(n151) );
  OAI2BB2XL U1075 ( .B0(n2110), .B1(n2241), .A0N(\register[3][6] ), .A1N(n2244), .Y(n152) );
  OAI2BB2XL U1076 ( .B0(n2107), .B1(n2241), .A0N(\register[3][7] ), .A1N(n2244), .Y(n153) );
  OAI2BB2XL U1077 ( .B0(n2104), .B1(n2242), .A0N(\register[3][8] ), .A1N(n2244), .Y(n154) );
  OAI2BB2XL U1078 ( .B0(n2101), .B1(n2242), .A0N(\register[3][9] ), .A1N(n2244), .Y(n155) );
  OAI2BB2XL U1079 ( .B0(n2098), .B1(n2242), .A0N(\register[3][10] ), .A1N(
        n2244), .Y(n156) );
  OAI2BB2XL U1080 ( .B0(n2095), .B1(n2242), .A0N(\register[3][11] ), .A1N(
        n2244), .Y(n157) );
  OAI2BB2XL U1081 ( .B0(n2092), .B1(n2242), .A0N(\register[3][12] ), .A1N(
        n2244), .Y(n158) );
  OAI2BB2XL U1082 ( .B0(n2089), .B1(n2242), .A0N(\register[3][13] ), .A1N(
        n2244), .Y(n159) );
  OAI2BB2XL U1083 ( .B0(n2086), .B1(n2242), .A0N(\register[3][14] ), .A1N(
        n2244), .Y(n160) );
  OAI2BB2XL U1084 ( .B0(n2083), .B1(n2242), .A0N(\register[3][15] ), .A1N(
        n2244), .Y(n161) );
  OAI2BB2XL U1085 ( .B0(n2080), .B1(n2243), .A0N(\register[3][16] ), .A1N(
        n2244), .Y(n162) );
  OAI2BB2XL U1086 ( .B0(n2077), .B1(n2243), .A0N(\register[3][17] ), .A1N(
        n2244), .Y(n163) );
  OAI2BB2XL U1087 ( .B0(n2074), .B1(n2242), .A0N(\register[3][18] ), .A1N(
        n2244), .Y(n164) );
  OAI2BB2XL U1088 ( .B0(n2071), .B1(n2243), .A0N(\register[3][19] ), .A1N(
        n2244), .Y(n165) );
  OAI2BB2XL U1089 ( .B0(n2068), .B1(n2243), .A0N(\register[3][20] ), .A1N(
        n2244), .Y(n166) );
  OAI2BB2XL U1090 ( .B0(n2065), .B1(n2243), .A0N(\register[3][21] ), .A1N(
        n2243), .Y(n167) );
  OAI2BB2XL U1091 ( .B0(n2062), .B1(n2243), .A0N(\register[3][22] ), .A1N(
        n2243), .Y(n168) );
  OAI2BB2XL U1092 ( .B0(n2059), .B1(n2243), .A0N(\register[3][23] ), .A1N(
        n2243), .Y(n169) );
  OAI2BB2XL U1093 ( .B0(n2056), .B1(n2243), .A0N(\register[3][24] ), .A1N(
        n2243), .Y(n170) );
  OAI2BB2XL U1094 ( .B0(n2053), .B1(n2242), .A0N(\register[3][25] ), .A1N(
        n2243), .Y(n171) );
  OAI2BB2XL U1095 ( .B0(n2050), .B1(n2242), .A0N(\register[3][26] ), .A1N(
        n2243), .Y(n172) );
  OAI2BB2XL U1096 ( .B0(n2047), .B1(n2242), .A0N(\register[3][27] ), .A1N(
        n2243), .Y(n173) );
  OAI2BB2XL U1097 ( .B0(n2044), .B1(n2241), .A0N(\register[3][28] ), .A1N(
        n2243), .Y(n174) );
  OAI2BB2XL U1098 ( .B0(n2041), .B1(n2241), .A0N(\register[3][29] ), .A1N(
        n2243), .Y(n175) );
  OAI2BB2XL U1099 ( .B0(n2038), .B1(n2241), .A0N(\register[3][30] ), .A1N(
        n2243), .Y(n176) );
  OAI2BB2XL U1100 ( .B0(n2035), .B1(n2241), .A0N(\register[3][31] ), .A1N(
        n2243), .Y(n177) );
  OAI2BB2XL U1101 ( .B0(n2128), .B1(n2237), .A0N(\register[4][0] ), .A1N(n2239), .Y(n178) );
  OAI2BB2XL U1102 ( .B0(n2125), .B1(n2237), .A0N(\register[4][1] ), .A1N(n2240), .Y(n179) );
  OAI2BB2XL U1103 ( .B0(n2122), .B1(n2237), .A0N(\register[4][2] ), .A1N(n2240), .Y(n180) );
  OAI2BB2XL U1104 ( .B0(n2119), .B1(n2237), .A0N(\register[4][3] ), .A1N(n2240), .Y(n181) );
  OAI2BB2XL U1105 ( .B0(n2116), .B1(n2237), .A0N(\register[4][4] ), .A1N(n2240), .Y(n182) );
  OAI2BB2XL U1106 ( .B0(n2113), .B1(n2237), .A0N(\register[4][5] ), .A1N(n2240), .Y(n183) );
  OAI2BB2XL U1107 ( .B0(n2110), .B1(n2237), .A0N(\register[4][6] ), .A1N(n2240), .Y(n184) );
  OAI2BB2XL U1108 ( .B0(n2107), .B1(n2237), .A0N(\register[4][7] ), .A1N(n2240), .Y(n185) );
  OAI2BB2XL U1109 ( .B0(n2104), .B1(n2238), .A0N(\register[4][8] ), .A1N(n2240), .Y(n186) );
  OAI2BB2XL U1110 ( .B0(n2101), .B1(n2238), .A0N(\register[4][9] ), .A1N(n2240), .Y(n187) );
  OAI2BB2XL U1111 ( .B0(n2098), .B1(n2238), .A0N(\register[4][10] ), .A1N(
        n2240), .Y(n188) );
  OAI2BB2XL U1112 ( .B0(n2095), .B1(n2238), .A0N(\register[4][11] ), .A1N(
        n2240), .Y(n189) );
  OAI2BB2XL U1113 ( .B0(n2092), .B1(n2238), .A0N(\register[4][12] ), .A1N(
        n2240), .Y(n190) );
  OAI2BB2XL U1114 ( .B0(n2089), .B1(n2238), .A0N(\register[4][13] ), .A1N(
        n2240), .Y(n191) );
  OAI2BB2XL U1115 ( .B0(n2086), .B1(n2238), .A0N(\register[4][14] ), .A1N(
        n2240), .Y(n192) );
  OAI2BB2XL U1116 ( .B0(n2083), .B1(n2238), .A0N(\register[4][15] ), .A1N(
        n2240), .Y(n193) );
  OAI2BB2XL U1117 ( .B0(n2080), .B1(n2239), .A0N(\register[4][16] ), .A1N(
        n2240), .Y(n194) );
  OAI2BB2XL U1118 ( .B0(n2077), .B1(n2239), .A0N(\register[4][17] ), .A1N(
        n2240), .Y(n195) );
  OAI2BB2XL U1119 ( .B0(n2074), .B1(n2238), .A0N(\register[4][18] ), .A1N(
        n2240), .Y(n196) );
  OAI2BB2XL U1120 ( .B0(n2071), .B1(n2239), .A0N(\register[4][19] ), .A1N(
        n2240), .Y(n197) );
  OAI2BB2XL U1121 ( .B0(n2068), .B1(n2239), .A0N(\register[4][20] ), .A1N(
        n2240), .Y(n198) );
  OAI2BB2XL U1122 ( .B0(n2065), .B1(n2239), .A0N(\register[4][21] ), .A1N(
        n2239), .Y(n199) );
  OAI2BB2XL U1123 ( .B0(n2062), .B1(n2239), .A0N(\register[4][22] ), .A1N(
        n2239), .Y(n200) );
  OAI2BB2XL U1124 ( .B0(n2059), .B1(n2239), .A0N(\register[4][23] ), .A1N(
        n2239), .Y(n201) );
  OAI2BB2XL U1125 ( .B0(n2056), .B1(n2239), .A0N(\register[4][24] ), .A1N(
        n2239), .Y(n202) );
  OAI2BB2XL U1126 ( .B0(n2053), .B1(n2238), .A0N(\register[4][25] ), .A1N(
        n2239), .Y(n203) );
  OAI2BB2XL U1127 ( .B0(n2050), .B1(n2238), .A0N(\register[4][26] ), .A1N(
        n2239), .Y(n204) );
  OAI2BB2XL U1128 ( .B0(n2047), .B1(n2238), .A0N(\register[4][27] ), .A1N(
        n2239), .Y(n205) );
  OAI2BB2XL U1129 ( .B0(n2044), .B1(n2237), .A0N(\register[4][28] ), .A1N(
        n2239), .Y(n206) );
  OAI2BB2XL U1130 ( .B0(n2041), .B1(n2237), .A0N(\register[4][29] ), .A1N(
        n2239), .Y(n207) );
  OAI2BB2XL U1131 ( .B0(n2038), .B1(n2237), .A0N(\register[4][30] ), .A1N(
        n2239), .Y(n208) );
  OAI2BB2XL U1132 ( .B0(n2035), .B1(n2237), .A0N(\register[4][31] ), .A1N(
        n2239), .Y(n209) );
  OAI2BB2XL U1133 ( .B0(n2128), .B1(n2233), .A0N(\register[5][0] ), .A1N(n2235), .Y(n210) );
  OAI2BB2XL U1134 ( .B0(n2125), .B1(n2233), .A0N(\register[5][1] ), .A1N(n2236), .Y(n211) );
  OAI2BB2XL U1135 ( .B0(n2122), .B1(n2233), .A0N(\register[5][2] ), .A1N(n2236), .Y(n212) );
  OAI2BB2XL U1136 ( .B0(n2119), .B1(n2233), .A0N(\register[5][3] ), .A1N(n2236), .Y(n213) );
  OAI2BB2XL U1137 ( .B0(n2116), .B1(n2233), .A0N(\register[5][4] ), .A1N(n2236), .Y(n214) );
  OAI2BB2XL U1138 ( .B0(n2113), .B1(n2233), .A0N(\register[5][5] ), .A1N(n2236), .Y(n215) );
  OAI2BB2XL U1139 ( .B0(n2110), .B1(n2233), .A0N(\register[5][6] ), .A1N(n2236), .Y(n216) );
  OAI2BB2XL U1140 ( .B0(n2107), .B1(n2233), .A0N(\register[5][7] ), .A1N(n2236), .Y(n217) );
  OAI2BB2XL U1141 ( .B0(n2104), .B1(n2234), .A0N(\register[5][8] ), .A1N(n2236), .Y(n218) );
  OAI2BB2XL U1142 ( .B0(n2101), .B1(n2234), .A0N(\register[5][9] ), .A1N(n2236), .Y(n219) );
  OAI2BB2XL U1143 ( .B0(n2098), .B1(n2234), .A0N(\register[5][10] ), .A1N(
        n2236), .Y(n220) );
  OAI2BB2XL U1144 ( .B0(n2095), .B1(n2234), .A0N(\register[5][11] ), .A1N(
        n2236), .Y(n221) );
  OAI2BB2XL U1145 ( .B0(n2092), .B1(n2234), .A0N(\register[5][12] ), .A1N(
        n2236), .Y(n222) );
  OAI2BB2XL U1146 ( .B0(n2089), .B1(n2234), .A0N(\register[5][13] ), .A1N(
        n2236), .Y(n223) );
  OAI2BB2XL U1147 ( .B0(n2086), .B1(n2234), .A0N(\register[5][14] ), .A1N(
        n2236), .Y(n224) );
  OAI2BB2XL U1148 ( .B0(n2083), .B1(n2234), .A0N(\register[5][15] ), .A1N(
        n2236), .Y(n225) );
  OAI2BB2XL U1149 ( .B0(n2080), .B1(n2235), .A0N(\register[5][16] ), .A1N(
        n2236), .Y(n226) );
  OAI2BB2XL U1150 ( .B0(n2077), .B1(n2235), .A0N(\register[5][17] ), .A1N(
        n2236), .Y(n227) );
  OAI2BB2XL U1151 ( .B0(n2074), .B1(n2234), .A0N(\register[5][18] ), .A1N(
        n2236), .Y(n228) );
  OAI2BB2XL U1152 ( .B0(n2071), .B1(n2235), .A0N(\register[5][19] ), .A1N(
        n2236), .Y(n229) );
  OAI2BB2XL U1153 ( .B0(n2068), .B1(n2235), .A0N(\register[5][20] ), .A1N(
        n2236), .Y(n230) );
  OAI2BB2XL U1154 ( .B0(n2065), .B1(n2235), .A0N(\register[5][21] ), .A1N(
        n2235), .Y(n231) );
  OAI2BB2XL U1155 ( .B0(n2062), .B1(n2235), .A0N(\register[5][22] ), .A1N(
        n2235), .Y(n232) );
  OAI2BB2XL U1156 ( .B0(n2059), .B1(n2235), .A0N(\register[5][23] ), .A1N(
        n2235), .Y(n233) );
  OAI2BB2XL U1157 ( .B0(n2056), .B1(n2235), .A0N(\register[5][24] ), .A1N(
        n2235), .Y(n234) );
  OAI2BB2XL U1158 ( .B0(n2053), .B1(n2234), .A0N(\register[5][25] ), .A1N(
        n2235), .Y(n235) );
  OAI2BB2XL U1159 ( .B0(n2050), .B1(n2234), .A0N(\register[5][26] ), .A1N(
        n2235), .Y(n236) );
  OAI2BB2XL U1160 ( .B0(n2047), .B1(n2234), .A0N(\register[5][27] ), .A1N(
        n2235), .Y(n237) );
  OAI2BB2XL U1161 ( .B0(n2044), .B1(n2233), .A0N(\register[5][28] ), .A1N(
        n2235), .Y(n238) );
  OAI2BB2XL U1162 ( .B0(n2041), .B1(n2233), .A0N(\register[5][29] ), .A1N(
        n2235), .Y(n239) );
  OAI2BB2XL U1163 ( .B0(n2038), .B1(n2233), .A0N(\register[5][30] ), .A1N(
        n2235), .Y(n240) );
  OAI2BB2XL U1164 ( .B0(n2035), .B1(n2233), .A0N(\register[5][31] ), .A1N(
        n2235), .Y(n241) );
  OAI2BB2XL U1165 ( .B0(n2128), .B1(n2229), .A0N(\register[6][0] ), .A1N(n2231), .Y(n242) );
  OAI2BB2XL U1166 ( .B0(n2125), .B1(n2229), .A0N(\register[6][1] ), .A1N(n2232), .Y(n243) );
  OAI2BB2XL U1167 ( .B0(n2122), .B1(n2229), .A0N(\register[6][2] ), .A1N(n2232), .Y(n244) );
  OAI2BB2XL U1168 ( .B0(n2119), .B1(n2229), .A0N(\register[6][3] ), .A1N(n2232), .Y(n245) );
  OAI2BB2XL U1169 ( .B0(n2116), .B1(n2229), .A0N(\register[6][4] ), .A1N(n2232), .Y(n246) );
  OAI2BB2XL U1170 ( .B0(n2113), .B1(n2229), .A0N(\register[6][5] ), .A1N(n2232), .Y(n247) );
  OAI2BB2XL U1171 ( .B0(n2110), .B1(n2229), .A0N(\register[6][6] ), .A1N(n2232), .Y(n248) );
  OAI2BB2XL U1172 ( .B0(n2107), .B1(n2229), .A0N(\register[6][7] ), .A1N(n2232), .Y(n249) );
  OAI2BB2XL U1173 ( .B0(n2104), .B1(n2230), .A0N(\register[6][8] ), .A1N(n2232), .Y(n250) );
  OAI2BB2XL U1174 ( .B0(n2101), .B1(n2230), .A0N(\register[6][9] ), .A1N(n2232), .Y(n251) );
  OAI2BB2XL U1175 ( .B0(n2098), .B1(n2230), .A0N(\register[6][10] ), .A1N(
        n2232), .Y(n252) );
  OAI2BB2XL U1176 ( .B0(n2095), .B1(n2230), .A0N(\register[6][11] ), .A1N(
        n2232), .Y(n253) );
  OAI2BB2XL U1177 ( .B0(n2092), .B1(n2230), .A0N(\register[6][12] ), .A1N(
        n2232), .Y(n254) );
  OAI2BB2XL U1178 ( .B0(n2089), .B1(n2230), .A0N(\register[6][13] ), .A1N(
        n2232), .Y(n255) );
  OAI2BB2XL U1179 ( .B0(n2086), .B1(n2230), .A0N(\register[6][14] ), .A1N(
        n2232), .Y(n256) );
  OAI2BB2XL U1180 ( .B0(n2083), .B1(n2230), .A0N(\register[6][15] ), .A1N(
        n2232), .Y(n257) );
  OAI2BB2XL U1181 ( .B0(n2080), .B1(n2231), .A0N(\register[6][16] ), .A1N(
        n2232), .Y(n258) );
  OAI2BB2XL U1182 ( .B0(n2077), .B1(n2231), .A0N(\register[6][17] ), .A1N(
        n2232), .Y(n259) );
  OAI2BB2XL U1183 ( .B0(n2074), .B1(n2230), .A0N(\register[6][18] ), .A1N(
        n2232), .Y(n260) );
  OAI2BB2XL U1184 ( .B0(n2071), .B1(n2231), .A0N(\register[6][19] ), .A1N(
        n2232), .Y(n261) );
  OAI2BB2XL U1185 ( .B0(n2068), .B1(n2231), .A0N(\register[6][20] ), .A1N(
        n2232), .Y(n262) );
  OAI2BB2XL U1186 ( .B0(n2065), .B1(n2231), .A0N(\register[6][21] ), .A1N(
        n2231), .Y(n263) );
  OAI2BB2XL U1187 ( .B0(n2062), .B1(n2231), .A0N(\register[6][22] ), .A1N(
        n2231), .Y(n264) );
  OAI2BB2XL U1188 ( .B0(n2059), .B1(n2231), .A0N(\register[6][23] ), .A1N(
        n2231), .Y(n265) );
  OAI2BB2XL U1189 ( .B0(n2056), .B1(n2231), .A0N(\register[6][24] ), .A1N(
        n2231), .Y(n266) );
  OAI2BB2XL U1190 ( .B0(n2053), .B1(n2230), .A0N(\register[6][25] ), .A1N(
        n2231), .Y(n267) );
  OAI2BB2XL U1191 ( .B0(n2050), .B1(n2230), .A0N(\register[6][26] ), .A1N(
        n2231), .Y(n268) );
  OAI2BB2XL U1192 ( .B0(n2047), .B1(n2230), .A0N(\register[6][27] ), .A1N(
        n2231), .Y(n269) );
  OAI2BB2XL U1193 ( .B0(n2044), .B1(n2229), .A0N(\register[6][28] ), .A1N(
        n2231), .Y(n270) );
  OAI2BB2XL U1194 ( .B0(n2041), .B1(n2229), .A0N(\register[6][29] ), .A1N(
        n2231), .Y(n271) );
  OAI2BB2XL U1195 ( .B0(n2038), .B1(n2229), .A0N(\register[6][30] ), .A1N(
        n2231), .Y(n272) );
  OAI2BB2XL U1196 ( .B0(n2035), .B1(n2229), .A0N(\register[6][31] ), .A1N(
        n2231), .Y(n273) );
  OAI2BB2XL U1197 ( .B0(n2128), .B1(n2225), .A0N(\register[7][0] ), .A1N(n2227), .Y(n274) );
  OAI2BB2XL U1198 ( .B0(n2125), .B1(n2225), .A0N(\register[7][1] ), .A1N(n2228), .Y(n275) );
  OAI2BB2XL U1199 ( .B0(n2122), .B1(n2225), .A0N(\register[7][2] ), .A1N(n2228), .Y(n276) );
  OAI2BB2XL U1200 ( .B0(n2119), .B1(n2225), .A0N(\register[7][3] ), .A1N(n2228), .Y(n277) );
  OAI2BB2XL U1201 ( .B0(n2116), .B1(n2225), .A0N(\register[7][4] ), .A1N(n2228), .Y(n278) );
  OAI2BB2XL U1202 ( .B0(n2113), .B1(n2225), .A0N(\register[7][5] ), .A1N(n2228), .Y(n279) );
  OAI2BB2XL U1203 ( .B0(n2110), .B1(n2225), .A0N(\register[7][6] ), .A1N(n2228), .Y(n280) );
  OAI2BB2XL U1204 ( .B0(n2107), .B1(n2225), .A0N(\register[7][7] ), .A1N(n2228), .Y(n281) );
  OAI2BB2XL U1205 ( .B0(n2104), .B1(n2226), .A0N(\register[7][8] ), .A1N(n2228), .Y(n282) );
  OAI2BB2XL U1206 ( .B0(n2101), .B1(n2226), .A0N(\register[7][9] ), .A1N(n2228), .Y(n283) );
  OAI2BB2XL U1207 ( .B0(n2098), .B1(n2226), .A0N(\register[7][10] ), .A1N(
        n2228), .Y(n284) );
  OAI2BB2XL U1208 ( .B0(n2095), .B1(n2226), .A0N(\register[7][11] ), .A1N(
        n2228), .Y(n285) );
  OAI2BB2XL U1209 ( .B0(n2092), .B1(n2226), .A0N(\register[7][12] ), .A1N(
        n2228), .Y(n286) );
  OAI2BB2XL U1210 ( .B0(n2089), .B1(n2226), .A0N(\register[7][13] ), .A1N(
        n2228), .Y(n287) );
  OAI2BB2XL U1211 ( .B0(n2086), .B1(n2226), .A0N(\register[7][14] ), .A1N(
        n2228), .Y(n288) );
  OAI2BB2XL U1212 ( .B0(n2083), .B1(n2226), .A0N(\register[7][15] ), .A1N(
        n2228), .Y(n289) );
  OAI2BB2XL U1213 ( .B0(n2080), .B1(n2227), .A0N(\register[7][16] ), .A1N(
        n2228), .Y(n290) );
  OAI2BB2XL U1214 ( .B0(n2077), .B1(n2227), .A0N(\register[7][17] ), .A1N(
        n2228), .Y(n291) );
  OAI2BB2XL U1215 ( .B0(n2074), .B1(n2226), .A0N(\register[7][18] ), .A1N(
        n2228), .Y(n292) );
  OAI2BB2XL U1216 ( .B0(n2071), .B1(n2227), .A0N(\register[7][19] ), .A1N(
        n2228), .Y(n293) );
  OAI2BB2XL U1217 ( .B0(n2068), .B1(n2227), .A0N(\register[7][20] ), .A1N(
        n2228), .Y(n294) );
  OAI2BB2XL U1218 ( .B0(n2065), .B1(n2227), .A0N(\register[7][21] ), .A1N(
        n2227), .Y(n295) );
  OAI2BB2XL U1219 ( .B0(n2062), .B1(n2227), .A0N(\register[7][22] ), .A1N(
        n2227), .Y(n296) );
  OAI2BB2XL U1220 ( .B0(n2059), .B1(n2227), .A0N(\register[7][23] ), .A1N(
        n2227), .Y(n297) );
  OAI2BB2XL U1221 ( .B0(n2056), .B1(n2227), .A0N(\register[7][24] ), .A1N(
        n2227), .Y(n298) );
  OAI2BB2XL U1222 ( .B0(n2053), .B1(n2226), .A0N(\register[7][25] ), .A1N(
        n2227), .Y(n299) );
  OAI2BB2XL U1223 ( .B0(n2050), .B1(n2226), .A0N(\register[7][26] ), .A1N(
        n2227), .Y(n300) );
  OAI2BB2XL U1224 ( .B0(n2047), .B1(n2226), .A0N(\register[7][27] ), .A1N(
        n2227), .Y(n301) );
  OAI2BB2XL U1225 ( .B0(n2044), .B1(n2225), .A0N(\register[7][28] ), .A1N(
        n2227), .Y(n302) );
  OAI2BB2XL U1226 ( .B0(n2041), .B1(n2225), .A0N(\register[7][29] ), .A1N(
        n2227), .Y(n303) );
  OAI2BB2XL U1227 ( .B0(n2038), .B1(n2225), .A0N(\register[7][30] ), .A1N(
        n2227), .Y(n304) );
  OAI2BB2XL U1228 ( .B0(n2035), .B1(n2225), .A0N(\register[7][31] ), .A1N(
        n2227), .Y(n305) );
  OAI2BB2XL U1229 ( .B0(n2127), .B1(n2221), .A0N(\register[8][0] ), .A1N(n2223), .Y(n306) );
  OAI2BB2XL U1230 ( .B0(n2124), .B1(n2221), .A0N(\register[8][1] ), .A1N(n2224), .Y(n307) );
  OAI2BB2XL U1231 ( .B0(n2121), .B1(n2221), .A0N(\register[8][2] ), .A1N(n2224), .Y(n308) );
  OAI2BB2XL U1232 ( .B0(n2118), .B1(n2221), .A0N(\register[8][3] ), .A1N(n2224), .Y(n309) );
  OAI2BB2XL U1233 ( .B0(n2115), .B1(n2221), .A0N(\register[8][4] ), .A1N(n2224), .Y(n310) );
  OAI2BB2XL U1234 ( .B0(n2112), .B1(n2221), .A0N(\register[8][5] ), .A1N(n2224), .Y(n311) );
  OAI2BB2XL U1235 ( .B0(n2109), .B1(n2221), .A0N(\register[8][6] ), .A1N(n2224), .Y(n312) );
  OAI2BB2XL U1236 ( .B0(n2106), .B1(n2221), .A0N(\register[8][7] ), .A1N(n2224), .Y(n313) );
  OAI2BB2XL U1237 ( .B0(n2103), .B1(n2222), .A0N(\register[8][8] ), .A1N(n2224), .Y(n314) );
  OAI2BB2XL U1238 ( .B0(n2100), .B1(n2222), .A0N(\register[8][9] ), .A1N(n2224), .Y(n315) );
  OAI2BB2XL U1239 ( .B0(n2097), .B1(n2222), .A0N(\register[8][10] ), .A1N(
        n2224), .Y(n316) );
  OAI2BB2XL U1240 ( .B0(n2094), .B1(n2222), .A0N(\register[8][11] ), .A1N(
        n2224), .Y(n317) );
  OAI2BB2XL U1241 ( .B0(n2091), .B1(n2222), .A0N(\register[8][12] ), .A1N(
        n2224), .Y(n318) );
  OAI2BB2XL U1242 ( .B0(n2088), .B1(n2222), .A0N(\register[8][13] ), .A1N(
        n2224), .Y(n319) );
  OAI2BB2XL U1243 ( .B0(n2085), .B1(n2222), .A0N(\register[8][14] ), .A1N(
        n2224), .Y(n320) );
  OAI2BB2XL U1244 ( .B0(n2082), .B1(n2222), .A0N(\register[8][15] ), .A1N(
        n2224), .Y(n321) );
  OAI2BB2XL U1245 ( .B0(n2079), .B1(n2223), .A0N(\register[8][16] ), .A1N(
        n2224), .Y(n322) );
  OAI2BB2XL U1246 ( .B0(n2076), .B1(n2223), .A0N(\register[8][17] ), .A1N(
        n2224), .Y(n323) );
  OAI2BB2XL U1247 ( .B0(n2073), .B1(n2222), .A0N(\register[8][18] ), .A1N(
        n2224), .Y(n324) );
  OAI2BB2XL U1248 ( .B0(n2070), .B1(n2223), .A0N(\register[8][19] ), .A1N(
        n2224), .Y(n325) );
  OAI2BB2XL U1249 ( .B0(n2067), .B1(n2223), .A0N(\register[8][20] ), .A1N(
        n2224), .Y(n326) );
  OAI2BB2XL U1250 ( .B0(n2064), .B1(n2223), .A0N(\register[8][21] ), .A1N(
        n2223), .Y(n327) );
  OAI2BB2XL U1251 ( .B0(n2061), .B1(n2223), .A0N(\register[8][22] ), .A1N(
        n2223), .Y(n328) );
  OAI2BB2XL U1252 ( .B0(n2058), .B1(n2223), .A0N(\register[8][23] ), .A1N(
        n2223), .Y(n329) );
  OAI2BB2XL U1253 ( .B0(n2055), .B1(n2223), .A0N(\register[8][24] ), .A1N(
        n2223), .Y(n330) );
  OAI2BB2XL U1254 ( .B0(n2052), .B1(n2222), .A0N(\register[8][25] ), .A1N(
        n2223), .Y(n331) );
  OAI2BB2XL U1255 ( .B0(n2049), .B1(n2222), .A0N(\register[8][26] ), .A1N(
        n2223), .Y(n332) );
  OAI2BB2XL U1256 ( .B0(n2046), .B1(n2222), .A0N(\register[8][27] ), .A1N(
        n2223), .Y(n333) );
  OAI2BB2XL U1257 ( .B0(n2043), .B1(n2221), .A0N(\register[8][28] ), .A1N(
        n2223), .Y(n334) );
  OAI2BB2XL U1258 ( .B0(n2040), .B1(n2221), .A0N(\register[8][29] ), .A1N(
        n2223), .Y(n335) );
  OAI2BB2XL U1259 ( .B0(n2037), .B1(n2221), .A0N(\register[8][30] ), .A1N(
        n2223), .Y(n336) );
  OAI2BB2XL U1260 ( .B0(n2034), .B1(n2221), .A0N(\register[8][31] ), .A1N(
        n2223), .Y(n337) );
  OAI2BB2XL U1261 ( .B0(n2127), .B1(n2217), .A0N(\register[9][0] ), .A1N(n2219), .Y(n338) );
  OAI2BB2XL U1262 ( .B0(n2124), .B1(n2217), .A0N(\register[9][1] ), .A1N(n2220), .Y(n339) );
  OAI2BB2XL U1263 ( .B0(n2121), .B1(n2217), .A0N(\register[9][2] ), .A1N(n2220), .Y(n340) );
  OAI2BB2XL U1264 ( .B0(n2118), .B1(n2217), .A0N(\register[9][3] ), .A1N(n2220), .Y(n341) );
  OAI2BB2XL U1265 ( .B0(n2115), .B1(n2217), .A0N(\register[9][4] ), .A1N(n2220), .Y(n342) );
  OAI2BB2XL U1266 ( .B0(n2112), .B1(n2217), .A0N(\register[9][5] ), .A1N(n2220), .Y(n343) );
  OAI2BB2XL U1267 ( .B0(n2109), .B1(n2217), .A0N(\register[9][6] ), .A1N(n2220), .Y(n344) );
  OAI2BB2XL U1268 ( .B0(n2106), .B1(n2217), .A0N(\register[9][7] ), .A1N(n2220), .Y(n345) );
  OAI2BB2XL U1269 ( .B0(n2103), .B1(n2218), .A0N(\register[9][8] ), .A1N(n2220), .Y(n346) );
  OAI2BB2XL U1270 ( .B0(n2100), .B1(n2218), .A0N(\register[9][9] ), .A1N(n2220), .Y(n347) );
  OAI2BB2XL U1271 ( .B0(n2097), .B1(n2218), .A0N(\register[9][10] ), .A1N(
        n2220), .Y(n348) );
  OAI2BB2XL U1272 ( .B0(n2094), .B1(n2218), .A0N(\register[9][11] ), .A1N(
        n2220), .Y(n349) );
  OAI2BB2XL U1273 ( .B0(n2091), .B1(n2218), .A0N(\register[9][12] ), .A1N(
        n2220), .Y(n350) );
  OAI2BB2XL U1274 ( .B0(n2088), .B1(n2218), .A0N(\register[9][13] ), .A1N(
        n2220), .Y(n351) );
  OAI2BB2XL U1275 ( .B0(n2085), .B1(n2218), .A0N(\register[9][14] ), .A1N(
        n2220), .Y(n352) );
  OAI2BB2XL U1276 ( .B0(n2082), .B1(n2218), .A0N(\register[9][15] ), .A1N(
        n2220), .Y(n353) );
  OAI2BB2XL U1277 ( .B0(n2079), .B1(n2219), .A0N(\register[9][16] ), .A1N(
        n2220), .Y(n354) );
  OAI2BB2XL U1278 ( .B0(n2076), .B1(n2219), .A0N(\register[9][17] ), .A1N(
        n2220), .Y(n355) );
  OAI2BB2XL U1279 ( .B0(n2073), .B1(n2218), .A0N(\register[9][18] ), .A1N(
        n2220), .Y(n356) );
  OAI2BB2XL U1280 ( .B0(n2070), .B1(n2219), .A0N(\register[9][19] ), .A1N(
        n2220), .Y(n357) );
  OAI2BB2XL U1281 ( .B0(n2067), .B1(n2219), .A0N(\register[9][20] ), .A1N(
        n2220), .Y(n358) );
  OAI2BB2XL U1282 ( .B0(n2064), .B1(n2219), .A0N(\register[9][21] ), .A1N(
        n2219), .Y(n359) );
  OAI2BB2XL U1283 ( .B0(n2061), .B1(n2219), .A0N(\register[9][22] ), .A1N(
        n2219), .Y(n360) );
  OAI2BB2XL U1284 ( .B0(n2058), .B1(n2219), .A0N(\register[9][23] ), .A1N(
        n2219), .Y(n361) );
  OAI2BB2XL U1285 ( .B0(n2055), .B1(n2219), .A0N(\register[9][24] ), .A1N(
        n2219), .Y(n362) );
  OAI2BB2XL U1286 ( .B0(n2052), .B1(n2218), .A0N(\register[9][25] ), .A1N(
        n2219), .Y(n363) );
  OAI2BB2XL U1287 ( .B0(n2049), .B1(n2218), .A0N(\register[9][26] ), .A1N(
        n2219), .Y(n364) );
  OAI2BB2XL U1288 ( .B0(n2046), .B1(n2218), .A0N(\register[9][27] ), .A1N(
        n2219), .Y(n365) );
  OAI2BB2XL U1289 ( .B0(n2043), .B1(n2217), .A0N(\register[9][28] ), .A1N(
        n2219), .Y(n366) );
  OAI2BB2XL U1290 ( .B0(n2040), .B1(n2217), .A0N(\register[9][29] ), .A1N(
        n2219), .Y(n367) );
  OAI2BB2XL U1291 ( .B0(n2037), .B1(n2217), .A0N(\register[9][30] ), .A1N(
        n2219), .Y(n368) );
  OAI2BB2XL U1292 ( .B0(n2034), .B1(n2217), .A0N(\register[9][31] ), .A1N(
        n2219), .Y(n369) );
  OAI2BB2XL U1293 ( .B0(n2127), .B1(n2213), .A0N(\register[10][0] ), .A1N(
        n2215), .Y(n370) );
  OAI2BB2XL U1294 ( .B0(n2124), .B1(n2213), .A0N(\register[10][1] ), .A1N(
        n2216), .Y(n371) );
  OAI2BB2XL U1295 ( .B0(n2121), .B1(n2213), .A0N(\register[10][2] ), .A1N(
        n2216), .Y(n372) );
  OAI2BB2XL U1296 ( .B0(n2118), .B1(n2213), .A0N(\register[10][3] ), .A1N(
        n2216), .Y(n373) );
  OAI2BB2XL U1297 ( .B0(n2115), .B1(n2213), .A0N(\register[10][4] ), .A1N(
        n2216), .Y(n374) );
  OAI2BB2XL U1298 ( .B0(n2112), .B1(n2213), .A0N(\register[10][5] ), .A1N(
        n2216), .Y(n375) );
  OAI2BB2XL U1299 ( .B0(n2109), .B1(n2213), .A0N(\register[10][6] ), .A1N(
        n2216), .Y(n376) );
  OAI2BB2XL U1300 ( .B0(n2106), .B1(n2213), .A0N(\register[10][7] ), .A1N(
        n2216), .Y(n377) );
  OAI2BB2XL U1301 ( .B0(n2103), .B1(n2214), .A0N(\register[10][8] ), .A1N(
        n2216), .Y(n378) );
  OAI2BB2XL U1302 ( .B0(n2100), .B1(n2214), .A0N(\register[10][9] ), .A1N(
        n2216), .Y(n379) );
  OAI2BB2XL U1303 ( .B0(n2097), .B1(n2214), .A0N(\register[10][10] ), .A1N(
        n2216), .Y(n380) );
  OAI2BB2XL U1304 ( .B0(n2094), .B1(n2214), .A0N(\register[10][11] ), .A1N(
        n2216), .Y(n381) );
  OAI2BB2XL U1305 ( .B0(n2091), .B1(n2214), .A0N(\register[10][12] ), .A1N(
        n2216), .Y(n382) );
  OAI2BB2XL U1306 ( .B0(n2088), .B1(n2214), .A0N(\register[10][13] ), .A1N(
        n2216), .Y(n383) );
  OAI2BB2XL U1307 ( .B0(n2085), .B1(n2214), .A0N(\register[10][14] ), .A1N(
        n2216), .Y(n384) );
  OAI2BB2XL U1308 ( .B0(n2082), .B1(n2214), .A0N(\register[10][15] ), .A1N(
        n2216), .Y(n385) );
  OAI2BB2XL U1309 ( .B0(n2079), .B1(n2215), .A0N(\register[10][16] ), .A1N(
        n2216), .Y(n386) );
  OAI2BB2XL U1310 ( .B0(n2076), .B1(n2215), .A0N(\register[10][17] ), .A1N(
        n2216), .Y(n387) );
  OAI2BB2XL U1311 ( .B0(n2073), .B1(n2214), .A0N(\register[10][18] ), .A1N(
        n2216), .Y(n388) );
  OAI2BB2XL U1312 ( .B0(n2070), .B1(n2215), .A0N(\register[10][19] ), .A1N(
        n2216), .Y(n389) );
  OAI2BB2XL U1313 ( .B0(n2067), .B1(n2215), .A0N(\register[10][20] ), .A1N(
        n2216), .Y(n390) );
  OAI2BB2XL U1314 ( .B0(n2064), .B1(n2215), .A0N(\register[10][21] ), .A1N(
        n2215), .Y(n391) );
  OAI2BB2XL U1315 ( .B0(n2061), .B1(n2215), .A0N(\register[10][22] ), .A1N(
        n2215), .Y(n392) );
  OAI2BB2XL U1316 ( .B0(n2058), .B1(n2215), .A0N(\register[10][23] ), .A1N(
        n2215), .Y(n393) );
  OAI2BB2XL U1317 ( .B0(n2055), .B1(n2215), .A0N(\register[10][24] ), .A1N(
        n2215), .Y(n394) );
  OAI2BB2XL U1318 ( .B0(n2052), .B1(n2214), .A0N(\register[10][25] ), .A1N(
        n2215), .Y(n395) );
  OAI2BB2XL U1319 ( .B0(n2049), .B1(n2214), .A0N(\register[10][26] ), .A1N(
        n2215), .Y(n396) );
  OAI2BB2XL U1320 ( .B0(n2046), .B1(n2214), .A0N(\register[10][27] ), .A1N(
        n2215), .Y(n397) );
  OAI2BB2XL U1321 ( .B0(n2043), .B1(n2213), .A0N(\register[10][28] ), .A1N(
        n2215), .Y(n398) );
  OAI2BB2XL U1322 ( .B0(n2040), .B1(n2213), .A0N(\register[10][29] ), .A1N(
        n2215), .Y(n399) );
  OAI2BB2XL U1323 ( .B0(n2037), .B1(n2213), .A0N(\register[10][30] ), .A1N(
        n2215), .Y(n400) );
  OAI2BB2XL U1324 ( .B0(n2034), .B1(n2213), .A0N(\register[10][31] ), .A1N(
        n2215), .Y(n401) );
  OAI2BB2XL U1325 ( .B0(n2127), .B1(n2209), .A0N(\register[11][0] ), .A1N(
        n2211), .Y(n402) );
  OAI2BB2XL U1326 ( .B0(n2124), .B1(n2209), .A0N(\register[11][1] ), .A1N(
        n2212), .Y(n403) );
  OAI2BB2XL U1327 ( .B0(n2121), .B1(n2209), .A0N(\register[11][2] ), .A1N(
        n2212), .Y(n404) );
  OAI2BB2XL U1328 ( .B0(n2118), .B1(n2209), .A0N(\register[11][3] ), .A1N(
        n2212), .Y(n405) );
  OAI2BB2XL U1329 ( .B0(n2115), .B1(n2209), .A0N(\register[11][4] ), .A1N(
        n2212), .Y(n406) );
  OAI2BB2XL U1330 ( .B0(n2112), .B1(n2209), .A0N(\register[11][5] ), .A1N(
        n2212), .Y(n407) );
  OAI2BB2XL U1331 ( .B0(n2109), .B1(n2209), .A0N(\register[11][6] ), .A1N(
        n2212), .Y(n408) );
  OAI2BB2XL U1332 ( .B0(n2106), .B1(n2209), .A0N(\register[11][7] ), .A1N(
        n2212), .Y(n409) );
  OAI2BB2XL U1333 ( .B0(n2103), .B1(n2210), .A0N(\register[11][8] ), .A1N(
        n2212), .Y(n410) );
  OAI2BB2XL U1334 ( .B0(n2100), .B1(n2210), .A0N(\register[11][9] ), .A1N(
        n2212), .Y(n411) );
  OAI2BB2XL U1335 ( .B0(n2097), .B1(n2210), .A0N(\register[11][10] ), .A1N(
        n2212), .Y(n412) );
  OAI2BB2XL U1336 ( .B0(n2094), .B1(n2210), .A0N(\register[11][11] ), .A1N(
        n2212), .Y(n413) );
  OAI2BB2XL U1337 ( .B0(n2091), .B1(n2210), .A0N(\register[11][12] ), .A1N(
        n2212), .Y(n414) );
  OAI2BB2XL U1338 ( .B0(n2088), .B1(n2210), .A0N(\register[11][13] ), .A1N(
        n2212), .Y(n415) );
  OAI2BB2XL U1339 ( .B0(n2085), .B1(n2210), .A0N(\register[11][14] ), .A1N(
        n2212), .Y(n416) );
  OAI2BB2XL U1340 ( .B0(n2082), .B1(n2210), .A0N(\register[11][15] ), .A1N(
        n2212), .Y(n417) );
  OAI2BB2XL U1341 ( .B0(n2079), .B1(n2211), .A0N(\register[11][16] ), .A1N(
        n2212), .Y(n418) );
  OAI2BB2XL U1342 ( .B0(n2076), .B1(n2211), .A0N(\register[11][17] ), .A1N(
        n2212), .Y(n419) );
  OAI2BB2XL U1343 ( .B0(n2073), .B1(n2210), .A0N(\register[11][18] ), .A1N(
        n2212), .Y(n420) );
  OAI2BB2XL U1344 ( .B0(n2070), .B1(n2211), .A0N(\register[11][19] ), .A1N(
        n2212), .Y(n421) );
  OAI2BB2XL U1345 ( .B0(n2067), .B1(n2211), .A0N(\register[11][20] ), .A1N(
        n2212), .Y(n422) );
  OAI2BB2XL U1346 ( .B0(n2064), .B1(n2211), .A0N(\register[11][21] ), .A1N(
        n2211), .Y(n423) );
  OAI2BB2XL U1347 ( .B0(n2061), .B1(n2211), .A0N(\register[11][22] ), .A1N(
        n2211), .Y(n424) );
  OAI2BB2XL U1348 ( .B0(n2058), .B1(n2211), .A0N(\register[11][23] ), .A1N(
        n2211), .Y(n425) );
  OAI2BB2XL U1349 ( .B0(n2055), .B1(n2211), .A0N(\register[11][24] ), .A1N(
        n2211), .Y(n426) );
  OAI2BB2XL U1350 ( .B0(n2052), .B1(n2210), .A0N(\register[11][25] ), .A1N(
        n2211), .Y(n427) );
  OAI2BB2XL U1351 ( .B0(n2049), .B1(n2210), .A0N(\register[11][26] ), .A1N(
        n2211), .Y(n428) );
  OAI2BB2XL U1352 ( .B0(n2046), .B1(n2210), .A0N(\register[11][27] ), .A1N(
        n2211), .Y(n429) );
  OAI2BB2XL U1353 ( .B0(n2043), .B1(n2209), .A0N(\register[11][28] ), .A1N(
        n2211), .Y(n430) );
  OAI2BB2XL U1354 ( .B0(n2040), .B1(n2209), .A0N(\register[11][29] ), .A1N(
        n2211), .Y(n431) );
  OAI2BB2XL U1355 ( .B0(n2037), .B1(n2209), .A0N(\register[11][30] ), .A1N(
        n2211), .Y(n432) );
  OAI2BB2XL U1356 ( .B0(n2034), .B1(n2209), .A0N(\register[11][31] ), .A1N(
        n2211), .Y(n433) );
  OAI2BB2XL U1357 ( .B0(n2127), .B1(n2205), .A0N(\register[12][0] ), .A1N(
        n2207), .Y(n434) );
  OAI2BB2XL U1358 ( .B0(n2124), .B1(n2205), .A0N(\register[12][1] ), .A1N(
        n2208), .Y(n435) );
  OAI2BB2XL U1359 ( .B0(n2121), .B1(n2205), .A0N(\register[12][2] ), .A1N(
        n2208), .Y(n436) );
  OAI2BB2XL U1360 ( .B0(n2118), .B1(n2205), .A0N(\register[12][3] ), .A1N(
        n2208), .Y(n437) );
  OAI2BB2XL U1361 ( .B0(n2115), .B1(n2205), .A0N(\register[12][4] ), .A1N(
        n2208), .Y(n438) );
  OAI2BB2XL U1362 ( .B0(n2112), .B1(n2205), .A0N(\register[12][5] ), .A1N(
        n2208), .Y(n439) );
  OAI2BB2XL U1363 ( .B0(n2109), .B1(n2205), .A0N(\register[12][6] ), .A1N(
        n2208), .Y(n440) );
  OAI2BB2XL U1364 ( .B0(n2106), .B1(n2205), .A0N(\register[12][7] ), .A1N(
        n2208), .Y(n441) );
  OAI2BB2XL U1365 ( .B0(n2103), .B1(n2206), .A0N(\register[12][8] ), .A1N(
        n2208), .Y(n442) );
  OAI2BB2XL U1366 ( .B0(n2100), .B1(n2206), .A0N(\register[12][9] ), .A1N(
        n2208), .Y(n443) );
  OAI2BB2XL U1367 ( .B0(n2097), .B1(n2206), .A0N(\register[12][10] ), .A1N(
        n2208), .Y(n444) );
  OAI2BB2XL U1368 ( .B0(n2094), .B1(n2206), .A0N(\register[12][11] ), .A1N(
        n2208), .Y(n445) );
  OAI2BB2XL U1369 ( .B0(n2091), .B1(n2206), .A0N(\register[12][12] ), .A1N(
        n2208), .Y(n446) );
  OAI2BB2XL U1370 ( .B0(n2088), .B1(n2206), .A0N(\register[12][13] ), .A1N(
        n2208), .Y(n447) );
  OAI2BB2XL U1371 ( .B0(n2085), .B1(n2206), .A0N(\register[12][14] ), .A1N(
        n2208), .Y(n448) );
  OAI2BB2XL U1372 ( .B0(n2082), .B1(n2206), .A0N(\register[12][15] ), .A1N(
        n2208), .Y(n449) );
  OAI2BB2XL U1373 ( .B0(n2079), .B1(n2207), .A0N(\register[12][16] ), .A1N(
        n2208), .Y(n450) );
  OAI2BB2XL U1374 ( .B0(n2076), .B1(n2207), .A0N(\register[12][17] ), .A1N(
        n2208), .Y(n451) );
  OAI2BB2XL U1375 ( .B0(n2073), .B1(n2206), .A0N(\register[12][18] ), .A1N(
        n2208), .Y(n452) );
  OAI2BB2XL U1376 ( .B0(n2070), .B1(n2207), .A0N(\register[12][19] ), .A1N(
        n2208), .Y(n453) );
  OAI2BB2XL U1377 ( .B0(n2067), .B1(n2207), .A0N(\register[12][20] ), .A1N(
        n2208), .Y(n454) );
  OAI2BB2XL U1378 ( .B0(n2064), .B1(n2207), .A0N(\register[12][21] ), .A1N(
        n2207), .Y(n455) );
  OAI2BB2XL U1379 ( .B0(n2061), .B1(n2207), .A0N(\register[12][22] ), .A1N(
        n2207), .Y(n456) );
  OAI2BB2XL U1380 ( .B0(n2058), .B1(n2207), .A0N(\register[12][23] ), .A1N(
        n2207), .Y(n457) );
  OAI2BB2XL U1381 ( .B0(n2055), .B1(n2207), .A0N(\register[12][24] ), .A1N(
        n2207), .Y(n458) );
  OAI2BB2XL U1382 ( .B0(n2052), .B1(n2206), .A0N(\register[12][25] ), .A1N(
        n2207), .Y(n459) );
  OAI2BB2XL U1383 ( .B0(n2049), .B1(n2206), .A0N(\register[12][26] ), .A1N(
        n2207), .Y(n460) );
  OAI2BB2XL U1384 ( .B0(n2046), .B1(n2206), .A0N(\register[12][27] ), .A1N(
        n2207), .Y(n461) );
  OAI2BB2XL U1385 ( .B0(n2043), .B1(n2205), .A0N(\register[12][28] ), .A1N(
        n2207), .Y(n462) );
  OAI2BB2XL U1386 ( .B0(n2040), .B1(n2205), .A0N(\register[12][29] ), .A1N(
        n2207), .Y(n463) );
  OAI2BB2XL U1387 ( .B0(n2037), .B1(n2205), .A0N(\register[12][30] ), .A1N(
        n2207), .Y(n464) );
  OAI2BB2XL U1388 ( .B0(n2034), .B1(n2205), .A0N(\register[12][31] ), .A1N(
        n2207), .Y(n465) );
  OAI2BB2XL U1389 ( .B0(n2127), .B1(n2201), .A0N(\register[13][0] ), .A1N(
        n2203), .Y(n466) );
  OAI2BB2XL U1390 ( .B0(n2124), .B1(n2201), .A0N(\register[13][1] ), .A1N(
        n2204), .Y(n467) );
  OAI2BB2XL U1391 ( .B0(n2121), .B1(n2201), .A0N(\register[13][2] ), .A1N(
        n2204), .Y(n468) );
  OAI2BB2XL U1392 ( .B0(n2118), .B1(n2201), .A0N(\register[13][3] ), .A1N(
        n2204), .Y(n469) );
  OAI2BB2XL U1393 ( .B0(n2115), .B1(n2201), .A0N(\register[13][4] ), .A1N(
        n2204), .Y(n470) );
  OAI2BB2XL U1394 ( .B0(n2112), .B1(n2201), .A0N(\register[13][5] ), .A1N(
        n2204), .Y(n471) );
  OAI2BB2XL U1395 ( .B0(n2109), .B1(n2201), .A0N(\register[13][6] ), .A1N(
        n2204), .Y(n472) );
  OAI2BB2XL U1396 ( .B0(n2106), .B1(n2201), .A0N(\register[13][7] ), .A1N(
        n2204), .Y(n473) );
  OAI2BB2XL U1397 ( .B0(n2103), .B1(n2202), .A0N(\register[13][8] ), .A1N(
        n2204), .Y(n474) );
  OAI2BB2XL U1398 ( .B0(n2100), .B1(n2202), .A0N(\register[13][9] ), .A1N(
        n2204), .Y(n475) );
  OAI2BB2XL U1399 ( .B0(n2097), .B1(n2202), .A0N(\register[13][10] ), .A1N(
        n2204), .Y(n476) );
  OAI2BB2XL U1400 ( .B0(n2094), .B1(n2202), .A0N(\register[13][11] ), .A1N(
        n2204), .Y(n477) );
  OAI2BB2XL U1401 ( .B0(n2091), .B1(n2202), .A0N(\register[13][12] ), .A1N(
        n2204), .Y(n478) );
  OAI2BB2XL U1402 ( .B0(n2088), .B1(n2202), .A0N(\register[13][13] ), .A1N(
        n2204), .Y(n479) );
  OAI2BB2XL U1403 ( .B0(n2085), .B1(n2202), .A0N(\register[13][14] ), .A1N(
        n2204), .Y(n480) );
  OAI2BB2XL U1404 ( .B0(n2082), .B1(n2202), .A0N(\register[13][15] ), .A1N(
        n2204), .Y(n481) );
  OAI2BB2XL U1405 ( .B0(n2079), .B1(n2203), .A0N(\register[13][16] ), .A1N(
        n2204), .Y(n482) );
  OAI2BB2XL U1406 ( .B0(n2076), .B1(n2203), .A0N(\register[13][17] ), .A1N(
        n2204), .Y(n483) );
  OAI2BB2XL U1407 ( .B0(n2073), .B1(n2202), .A0N(\register[13][18] ), .A1N(
        n2204), .Y(n484) );
  OAI2BB2XL U1408 ( .B0(n2070), .B1(n2203), .A0N(\register[13][19] ), .A1N(
        n2204), .Y(n485) );
  OAI2BB2XL U1409 ( .B0(n2067), .B1(n2203), .A0N(\register[13][20] ), .A1N(
        n2204), .Y(n486) );
  OAI2BB2XL U1410 ( .B0(n2064), .B1(n2203), .A0N(\register[13][21] ), .A1N(
        n2203), .Y(n487) );
  OAI2BB2XL U1411 ( .B0(n2061), .B1(n2203), .A0N(\register[13][22] ), .A1N(
        n2203), .Y(n488) );
  OAI2BB2XL U1412 ( .B0(n2058), .B1(n2203), .A0N(\register[13][23] ), .A1N(
        n2203), .Y(n489) );
  OAI2BB2XL U1413 ( .B0(n2055), .B1(n2203), .A0N(\register[13][24] ), .A1N(
        n2203), .Y(n490) );
  OAI2BB2XL U1414 ( .B0(n2052), .B1(n2202), .A0N(\register[13][25] ), .A1N(
        n2203), .Y(n491) );
  OAI2BB2XL U1415 ( .B0(n2049), .B1(n2202), .A0N(\register[13][26] ), .A1N(
        n2203), .Y(n492) );
  OAI2BB2XL U1416 ( .B0(n2046), .B1(n2202), .A0N(\register[13][27] ), .A1N(
        n2203), .Y(n493) );
  OAI2BB2XL U1417 ( .B0(n2043), .B1(n2201), .A0N(\register[13][28] ), .A1N(
        n2203), .Y(n494) );
  OAI2BB2XL U1418 ( .B0(n2040), .B1(n2201), .A0N(\register[13][29] ), .A1N(
        n2203), .Y(n495) );
  OAI2BB2XL U1419 ( .B0(n2037), .B1(n2201), .A0N(\register[13][30] ), .A1N(
        n2203), .Y(n496) );
  OAI2BB2XL U1420 ( .B0(n2034), .B1(n2201), .A0N(\register[13][31] ), .A1N(
        n2203), .Y(n497) );
  OAI2BB2XL U1421 ( .B0(n2127), .B1(n2197), .A0N(\register[14][0] ), .A1N(
        n2199), .Y(n498) );
  OAI2BB2XL U1422 ( .B0(n2124), .B1(n2197), .A0N(\register[14][1] ), .A1N(
        n2200), .Y(n499) );
  OAI2BB2XL U1423 ( .B0(n2121), .B1(n2197), .A0N(\register[14][2] ), .A1N(
        n2200), .Y(n500) );
  OAI2BB2XL U1424 ( .B0(n2118), .B1(n2197), .A0N(\register[14][3] ), .A1N(
        n2200), .Y(n501) );
  OAI2BB2XL U1425 ( .B0(n2115), .B1(n2197), .A0N(\register[14][4] ), .A1N(
        n2200), .Y(n502) );
  OAI2BB2XL U1426 ( .B0(n2112), .B1(n2197), .A0N(\register[14][5] ), .A1N(
        n2200), .Y(n503) );
  OAI2BB2XL U1427 ( .B0(n2109), .B1(n2197), .A0N(\register[14][6] ), .A1N(
        n2200), .Y(n504) );
  OAI2BB2XL U1428 ( .B0(n2106), .B1(n2197), .A0N(\register[14][7] ), .A1N(
        n2200), .Y(n505) );
  OAI2BB2XL U1429 ( .B0(n2103), .B1(n2198), .A0N(\register[14][8] ), .A1N(
        n2200), .Y(n506) );
  OAI2BB2XL U1430 ( .B0(n2100), .B1(n2198), .A0N(\register[14][9] ), .A1N(
        n2200), .Y(n507) );
  OAI2BB2XL U1431 ( .B0(n2097), .B1(n2198), .A0N(\register[14][10] ), .A1N(
        n2200), .Y(n508) );
  OAI2BB2XL U1432 ( .B0(n2094), .B1(n2198), .A0N(\register[14][11] ), .A1N(
        n2200), .Y(n509) );
  OAI2BB2XL U1433 ( .B0(n2091), .B1(n2198), .A0N(\register[14][12] ), .A1N(
        n2200), .Y(n510) );
  OAI2BB2XL U1434 ( .B0(n2088), .B1(n2198), .A0N(\register[14][13] ), .A1N(
        n2200), .Y(n511) );
  OAI2BB2XL U1435 ( .B0(n2085), .B1(n2198), .A0N(\register[14][14] ), .A1N(
        n2200), .Y(n512) );
  OAI2BB2XL U1436 ( .B0(n2082), .B1(n2198), .A0N(\register[14][15] ), .A1N(
        n2200), .Y(n513) );
  OAI2BB2XL U1437 ( .B0(n2079), .B1(n2199), .A0N(\register[14][16] ), .A1N(
        n2200), .Y(n514) );
  OAI2BB2XL U1438 ( .B0(n2076), .B1(n2199), .A0N(\register[14][17] ), .A1N(
        n2200), .Y(n515) );
  OAI2BB2XL U1439 ( .B0(n2073), .B1(n2198), .A0N(\register[14][18] ), .A1N(
        n2200), .Y(n516) );
  OAI2BB2XL U1440 ( .B0(n2070), .B1(n2199), .A0N(\register[14][19] ), .A1N(
        n2200), .Y(n517) );
  OAI2BB2XL U1441 ( .B0(n2067), .B1(n2199), .A0N(\register[14][20] ), .A1N(
        n2200), .Y(n518) );
  OAI2BB2XL U1442 ( .B0(n2064), .B1(n2199), .A0N(\register[14][21] ), .A1N(
        n2199), .Y(n519) );
  OAI2BB2XL U1443 ( .B0(n2061), .B1(n2199), .A0N(\register[14][22] ), .A1N(
        n2199), .Y(n520) );
  OAI2BB2XL U1444 ( .B0(n2058), .B1(n2199), .A0N(\register[14][23] ), .A1N(
        n2199), .Y(n521) );
  OAI2BB2XL U1445 ( .B0(n2055), .B1(n2199), .A0N(\register[14][24] ), .A1N(
        n2199), .Y(n522) );
  OAI2BB2XL U1446 ( .B0(n2052), .B1(n2198), .A0N(\register[14][25] ), .A1N(
        n2199), .Y(n523) );
  OAI2BB2XL U1447 ( .B0(n2049), .B1(n2198), .A0N(\register[14][26] ), .A1N(
        n2199), .Y(n524) );
  OAI2BB2XL U1448 ( .B0(n2046), .B1(n2198), .A0N(\register[14][27] ), .A1N(
        n2199), .Y(n525) );
  OAI2BB2XL U1449 ( .B0(n2043), .B1(n2197), .A0N(\register[14][28] ), .A1N(
        n2199), .Y(n526) );
  OAI2BB2XL U1450 ( .B0(n2040), .B1(n2197), .A0N(\register[14][29] ), .A1N(
        n2199), .Y(n527) );
  OAI2BB2XL U1451 ( .B0(n2037), .B1(n2197), .A0N(\register[14][30] ), .A1N(
        n2199), .Y(n528) );
  OAI2BB2XL U1452 ( .B0(n2034), .B1(n2197), .A0N(\register[14][31] ), .A1N(
        n2199), .Y(n529) );
  OAI2BB2XL U1453 ( .B0(n2127), .B1(n2193), .A0N(\register[15][0] ), .A1N(
        n2195), .Y(n530) );
  OAI2BB2XL U1454 ( .B0(n2124), .B1(n2193), .A0N(\register[15][1] ), .A1N(
        n2196), .Y(n531) );
  OAI2BB2XL U1455 ( .B0(n2121), .B1(n2193), .A0N(\register[15][2] ), .A1N(
        n2196), .Y(n532) );
  OAI2BB2XL U1456 ( .B0(n2118), .B1(n2193), .A0N(\register[15][3] ), .A1N(
        n2196), .Y(n533) );
  OAI2BB2XL U1457 ( .B0(n2115), .B1(n2193), .A0N(\register[15][4] ), .A1N(
        n2196), .Y(n534) );
  OAI2BB2XL U1458 ( .B0(n2112), .B1(n2193), .A0N(\register[15][5] ), .A1N(
        n2196), .Y(n535) );
  OAI2BB2XL U1459 ( .B0(n2109), .B1(n2193), .A0N(\register[15][6] ), .A1N(
        n2196), .Y(n536) );
  OAI2BB2XL U1460 ( .B0(n2106), .B1(n2193), .A0N(\register[15][7] ), .A1N(
        n2196), .Y(n537) );
  OAI2BB2XL U1461 ( .B0(n2103), .B1(n2194), .A0N(\register[15][8] ), .A1N(
        n2196), .Y(n538) );
  OAI2BB2XL U1462 ( .B0(n2100), .B1(n2194), .A0N(\register[15][9] ), .A1N(
        n2196), .Y(n539) );
  OAI2BB2XL U1463 ( .B0(n2097), .B1(n2194), .A0N(\register[15][10] ), .A1N(
        n2196), .Y(n540) );
  OAI2BB2XL U1464 ( .B0(n2094), .B1(n2194), .A0N(\register[15][11] ), .A1N(
        n2196), .Y(n541) );
  OAI2BB2XL U1465 ( .B0(n2091), .B1(n2194), .A0N(\register[15][12] ), .A1N(
        n2196), .Y(n542) );
  OAI2BB2XL U1466 ( .B0(n2088), .B1(n2194), .A0N(\register[15][13] ), .A1N(
        n2196), .Y(n543) );
  OAI2BB2XL U1467 ( .B0(n2085), .B1(n2194), .A0N(\register[15][14] ), .A1N(
        n2196), .Y(n544) );
  OAI2BB2XL U1468 ( .B0(n2082), .B1(n2194), .A0N(\register[15][15] ), .A1N(
        n2196), .Y(n545) );
  OAI2BB2XL U1469 ( .B0(n2079), .B1(n2195), .A0N(\register[15][16] ), .A1N(
        n2196), .Y(n546) );
  OAI2BB2XL U1470 ( .B0(n2076), .B1(n2195), .A0N(\register[15][17] ), .A1N(
        n2196), .Y(n547) );
  OAI2BB2XL U1471 ( .B0(n2073), .B1(n2194), .A0N(\register[15][18] ), .A1N(
        n2196), .Y(n548) );
  OAI2BB2XL U1472 ( .B0(n2070), .B1(n2195), .A0N(\register[15][19] ), .A1N(
        n2196), .Y(n549) );
  OAI2BB2XL U1473 ( .B0(n2067), .B1(n2195), .A0N(\register[15][20] ), .A1N(
        n2196), .Y(n550) );
  OAI2BB2XL U1474 ( .B0(n2064), .B1(n2195), .A0N(\register[15][21] ), .A1N(
        n2195), .Y(n551) );
  OAI2BB2XL U1475 ( .B0(n2061), .B1(n2195), .A0N(\register[15][22] ), .A1N(
        n2195), .Y(n552) );
  OAI2BB2XL U1476 ( .B0(n2058), .B1(n2195), .A0N(\register[15][23] ), .A1N(
        n2195), .Y(n553) );
  OAI2BB2XL U1477 ( .B0(n2055), .B1(n2195), .A0N(\register[15][24] ), .A1N(
        n2195), .Y(n554) );
  OAI2BB2XL U1478 ( .B0(n2052), .B1(n2194), .A0N(\register[15][25] ), .A1N(
        n2195), .Y(n555) );
  OAI2BB2XL U1479 ( .B0(n2049), .B1(n2194), .A0N(\register[15][26] ), .A1N(
        n2195), .Y(n556) );
  OAI2BB2XL U1480 ( .B0(n2046), .B1(n2194), .A0N(\register[15][27] ), .A1N(
        n2195), .Y(n557) );
  OAI2BB2XL U1481 ( .B0(n2043), .B1(n2193), .A0N(\register[15][28] ), .A1N(
        n2195), .Y(n558) );
  OAI2BB2XL U1482 ( .B0(n2040), .B1(n2193), .A0N(\register[15][29] ), .A1N(
        n2195), .Y(n559) );
  OAI2BB2XL U1483 ( .B0(n2037), .B1(n2193), .A0N(\register[15][30] ), .A1N(
        n2195), .Y(n560) );
  OAI2BB2XL U1484 ( .B0(n2034), .B1(n2193), .A0N(\register[15][31] ), .A1N(
        n2195), .Y(n561) );
  OAI2BB2XL U1485 ( .B0(n2127), .B1(n2189), .A0N(\register[16][0] ), .A1N(
        n2191), .Y(n562) );
  OAI2BB2XL U1486 ( .B0(n2124), .B1(n2189), .A0N(\register[16][1] ), .A1N(
        n2192), .Y(n563) );
  OAI2BB2XL U1487 ( .B0(n2121), .B1(n2189), .A0N(\register[16][2] ), .A1N(
        n2192), .Y(n564) );
  OAI2BB2XL U1488 ( .B0(n2118), .B1(n2189), .A0N(\register[16][3] ), .A1N(
        n2192), .Y(n565) );
  OAI2BB2XL U1489 ( .B0(n2115), .B1(n2189), .A0N(\register[16][4] ), .A1N(
        n2192), .Y(n566) );
  OAI2BB2XL U1490 ( .B0(n2112), .B1(n2189), .A0N(\register[16][5] ), .A1N(
        n2192), .Y(n567) );
  OAI2BB2XL U1491 ( .B0(n2109), .B1(n2189), .A0N(\register[16][6] ), .A1N(
        n2192), .Y(n568) );
  OAI2BB2XL U1492 ( .B0(n2106), .B1(n2189), .A0N(\register[16][7] ), .A1N(
        n2192), .Y(n569) );
  OAI2BB2XL U1493 ( .B0(n2103), .B1(n2190), .A0N(\register[16][8] ), .A1N(
        n2192), .Y(n570) );
  OAI2BB2XL U1494 ( .B0(n2100), .B1(n2190), .A0N(\register[16][9] ), .A1N(
        n2192), .Y(n571) );
  OAI2BB2XL U1495 ( .B0(n2097), .B1(n2190), .A0N(\register[16][10] ), .A1N(
        n2192), .Y(n572) );
  OAI2BB2XL U1496 ( .B0(n2094), .B1(n2190), .A0N(\register[16][11] ), .A1N(
        n2192), .Y(n573) );
  OAI2BB2XL U1497 ( .B0(n2091), .B1(n2190), .A0N(\register[16][12] ), .A1N(
        n2192), .Y(n574) );
  OAI2BB2XL U1498 ( .B0(n2088), .B1(n2190), .A0N(\register[16][13] ), .A1N(
        n2192), .Y(n575) );
  OAI2BB2XL U1499 ( .B0(n2085), .B1(n2190), .A0N(\register[16][14] ), .A1N(
        n2192), .Y(n576) );
  OAI2BB2XL U1500 ( .B0(n2082), .B1(n2190), .A0N(\register[16][15] ), .A1N(
        n2192), .Y(n577) );
  OAI2BB2XL U1501 ( .B0(n2079), .B1(n2191), .A0N(\register[16][16] ), .A1N(
        n2192), .Y(n578) );
  OAI2BB2XL U1502 ( .B0(n2076), .B1(n2191), .A0N(\register[16][17] ), .A1N(
        n2192), .Y(n579) );
  OAI2BB2XL U1503 ( .B0(n2073), .B1(n2190), .A0N(\register[16][18] ), .A1N(
        n2192), .Y(n580) );
  OAI2BB2XL U1504 ( .B0(n2070), .B1(n2191), .A0N(\register[16][19] ), .A1N(
        n2192), .Y(n581) );
  OAI2BB2XL U1505 ( .B0(n2067), .B1(n2191), .A0N(\register[16][20] ), .A1N(
        n2192), .Y(n582) );
  OAI2BB2XL U1506 ( .B0(n2064), .B1(n2191), .A0N(\register[16][21] ), .A1N(
        n2191), .Y(n583) );
  OAI2BB2XL U1507 ( .B0(n2061), .B1(n2191), .A0N(\register[16][22] ), .A1N(
        n2191), .Y(n584) );
  OAI2BB2XL U1508 ( .B0(n2058), .B1(n2191), .A0N(\register[16][23] ), .A1N(
        n2191), .Y(n585) );
  OAI2BB2XL U1509 ( .B0(n2055), .B1(n2191), .A0N(\register[16][24] ), .A1N(
        n2191), .Y(n586) );
  OAI2BB2XL U1510 ( .B0(n2052), .B1(n2190), .A0N(\register[16][25] ), .A1N(
        n2191), .Y(n587) );
  OAI2BB2XL U1511 ( .B0(n2049), .B1(n2190), .A0N(\register[16][26] ), .A1N(
        n2191), .Y(n588) );
  OAI2BB2XL U1512 ( .B0(n2046), .B1(n2190), .A0N(\register[16][27] ), .A1N(
        n2191), .Y(n589) );
  OAI2BB2XL U1513 ( .B0(n2043), .B1(n2189), .A0N(\register[16][28] ), .A1N(
        n2191), .Y(n590) );
  OAI2BB2XL U1514 ( .B0(n2040), .B1(n2189), .A0N(\register[16][29] ), .A1N(
        n2191), .Y(n591) );
  OAI2BB2XL U1515 ( .B0(n2037), .B1(n2189), .A0N(\register[16][30] ), .A1N(
        n2191), .Y(n592) );
  OAI2BB2XL U1516 ( .B0(n2034), .B1(n2189), .A0N(\register[16][31] ), .A1N(
        n2191), .Y(n593) );
  OAI2BB2XL U1517 ( .B0(n2127), .B1(n2185), .A0N(\register[17][0] ), .A1N(
        n2187), .Y(n594) );
  OAI2BB2XL U1518 ( .B0(n2124), .B1(n2185), .A0N(\register[17][1] ), .A1N(
        n2188), .Y(n595) );
  OAI2BB2XL U1519 ( .B0(n2121), .B1(n2185), .A0N(\register[17][2] ), .A1N(
        n2188), .Y(n596) );
  OAI2BB2XL U1520 ( .B0(n2118), .B1(n2185), .A0N(\register[17][3] ), .A1N(
        n2188), .Y(n597) );
  OAI2BB2XL U1521 ( .B0(n2115), .B1(n2185), .A0N(\register[17][4] ), .A1N(
        n2188), .Y(n598) );
  OAI2BB2XL U1522 ( .B0(n2112), .B1(n2185), .A0N(\register[17][5] ), .A1N(
        n2188), .Y(n599) );
  OAI2BB2XL U1523 ( .B0(n2109), .B1(n2185), .A0N(\register[17][6] ), .A1N(
        n2188), .Y(n600) );
  OAI2BB2XL U1524 ( .B0(n2106), .B1(n2185), .A0N(\register[17][7] ), .A1N(
        n2188), .Y(n601) );
  OAI2BB2XL U1525 ( .B0(n2103), .B1(n2186), .A0N(\register[17][8] ), .A1N(
        n2188), .Y(n602) );
  OAI2BB2XL U1526 ( .B0(n2100), .B1(n2186), .A0N(\register[17][9] ), .A1N(
        n2188), .Y(n603) );
  OAI2BB2XL U1527 ( .B0(n2097), .B1(n2186), .A0N(\register[17][10] ), .A1N(
        n2188), .Y(n604) );
  OAI2BB2XL U1528 ( .B0(n2094), .B1(n2186), .A0N(\register[17][11] ), .A1N(
        n2188), .Y(n605) );
  OAI2BB2XL U1529 ( .B0(n2091), .B1(n2186), .A0N(\register[17][12] ), .A1N(
        n2188), .Y(n606) );
  OAI2BB2XL U1530 ( .B0(n2088), .B1(n2186), .A0N(\register[17][13] ), .A1N(
        n2188), .Y(n607) );
  OAI2BB2XL U1531 ( .B0(n2085), .B1(n2186), .A0N(\register[17][14] ), .A1N(
        n2188), .Y(n608) );
  OAI2BB2XL U1532 ( .B0(n2082), .B1(n2186), .A0N(\register[17][15] ), .A1N(
        n2188), .Y(n609) );
  OAI2BB2XL U1533 ( .B0(n2079), .B1(n2187), .A0N(\register[17][16] ), .A1N(
        n2188), .Y(n610) );
  OAI2BB2XL U1534 ( .B0(n2076), .B1(n2187), .A0N(\register[17][17] ), .A1N(
        n2188), .Y(n611) );
  OAI2BB2XL U1535 ( .B0(n2073), .B1(n2186), .A0N(\register[17][18] ), .A1N(
        n2188), .Y(n612) );
  OAI2BB2XL U1536 ( .B0(n2070), .B1(n2187), .A0N(\register[17][19] ), .A1N(
        n2188), .Y(n613) );
  OAI2BB2XL U1537 ( .B0(n2067), .B1(n2187), .A0N(\register[17][20] ), .A1N(
        n2188), .Y(n614) );
  OAI2BB2XL U1538 ( .B0(n2064), .B1(n2187), .A0N(\register[17][21] ), .A1N(
        n2187), .Y(n615) );
  OAI2BB2XL U1539 ( .B0(n2061), .B1(n2187), .A0N(\register[17][22] ), .A1N(
        n2187), .Y(n616) );
  OAI2BB2XL U1540 ( .B0(n2058), .B1(n2187), .A0N(\register[17][23] ), .A1N(
        n2187), .Y(n617) );
  OAI2BB2XL U1541 ( .B0(n2055), .B1(n2187), .A0N(\register[17][24] ), .A1N(
        n2187), .Y(n618) );
  OAI2BB2XL U1542 ( .B0(n2052), .B1(n2186), .A0N(\register[17][25] ), .A1N(
        n2187), .Y(n619) );
  OAI2BB2XL U1543 ( .B0(n2049), .B1(n2186), .A0N(\register[17][26] ), .A1N(
        n2187), .Y(n620) );
  OAI2BB2XL U1544 ( .B0(n2046), .B1(n2186), .A0N(\register[17][27] ), .A1N(
        n2187), .Y(n621) );
  OAI2BB2XL U1545 ( .B0(n2043), .B1(n2185), .A0N(\register[17][28] ), .A1N(
        n2187), .Y(n622) );
  OAI2BB2XL U1546 ( .B0(n2040), .B1(n2185), .A0N(\register[17][29] ), .A1N(
        n2187), .Y(n623) );
  OAI2BB2XL U1547 ( .B0(n2037), .B1(n2185), .A0N(\register[17][30] ), .A1N(
        n2187), .Y(n624) );
  OAI2BB2XL U1548 ( .B0(n2034), .B1(n2185), .A0N(\register[17][31] ), .A1N(
        n2187), .Y(n625) );
  OAI2BB2XL U1549 ( .B0(n2127), .B1(n2181), .A0N(\register[18][0] ), .A1N(
        n2183), .Y(n626) );
  OAI2BB2XL U1550 ( .B0(n2124), .B1(n2181), .A0N(\register[18][1] ), .A1N(
        n2184), .Y(n627) );
  OAI2BB2XL U1551 ( .B0(n2121), .B1(n2181), .A0N(\register[18][2] ), .A1N(
        n2184), .Y(n628) );
  OAI2BB2XL U1552 ( .B0(n2118), .B1(n2181), .A0N(\register[18][3] ), .A1N(
        n2184), .Y(n629) );
  OAI2BB2XL U1553 ( .B0(n2115), .B1(n2181), .A0N(\register[18][4] ), .A1N(
        n2184), .Y(n630) );
  OAI2BB2XL U1554 ( .B0(n2112), .B1(n2181), .A0N(\register[18][5] ), .A1N(
        n2184), .Y(n631) );
  OAI2BB2XL U1555 ( .B0(n2109), .B1(n2181), .A0N(\register[18][6] ), .A1N(
        n2184), .Y(n632) );
  OAI2BB2XL U1556 ( .B0(n2106), .B1(n2181), .A0N(\register[18][7] ), .A1N(
        n2184), .Y(n633) );
  OAI2BB2XL U1557 ( .B0(n2103), .B1(n2182), .A0N(\register[18][8] ), .A1N(
        n2184), .Y(n634) );
  OAI2BB2XL U1558 ( .B0(n2100), .B1(n2182), .A0N(\register[18][9] ), .A1N(
        n2184), .Y(n635) );
  OAI2BB2XL U1559 ( .B0(n2097), .B1(n2182), .A0N(\register[18][10] ), .A1N(
        n2184), .Y(n636) );
  OAI2BB2XL U1560 ( .B0(n2094), .B1(n2182), .A0N(\register[18][11] ), .A1N(
        n2184), .Y(n637) );
  OAI2BB2XL U1561 ( .B0(n2091), .B1(n2182), .A0N(\register[18][12] ), .A1N(
        n2184), .Y(n638) );
  OAI2BB2XL U1562 ( .B0(n2088), .B1(n2182), .A0N(\register[18][13] ), .A1N(
        n2184), .Y(n639) );
  OAI2BB2XL U1563 ( .B0(n2085), .B1(n2182), .A0N(\register[18][14] ), .A1N(
        n2184), .Y(n640) );
  OAI2BB2XL U1564 ( .B0(n2082), .B1(n2182), .A0N(\register[18][15] ), .A1N(
        n2184), .Y(n641) );
  OAI2BB2XL U1565 ( .B0(n2079), .B1(n2183), .A0N(\register[18][16] ), .A1N(
        n2184), .Y(n642) );
  OAI2BB2XL U1566 ( .B0(n2076), .B1(n2183), .A0N(\register[18][17] ), .A1N(
        n2184), .Y(n643) );
  OAI2BB2XL U1567 ( .B0(n2073), .B1(n2182), .A0N(\register[18][18] ), .A1N(
        n2184), .Y(n644) );
  OAI2BB2XL U1568 ( .B0(n2070), .B1(n2183), .A0N(\register[18][19] ), .A1N(
        n2184), .Y(n645) );
  OAI2BB2XL U1569 ( .B0(n2067), .B1(n2183), .A0N(\register[18][20] ), .A1N(
        n2184), .Y(n646) );
  OAI2BB2XL U1570 ( .B0(n2064), .B1(n2183), .A0N(\register[18][21] ), .A1N(
        n2183), .Y(n647) );
  OAI2BB2XL U1571 ( .B0(n2061), .B1(n2183), .A0N(\register[18][22] ), .A1N(
        n2183), .Y(n648) );
  OAI2BB2XL U1572 ( .B0(n2058), .B1(n2183), .A0N(\register[18][23] ), .A1N(
        n2183), .Y(n649) );
  OAI2BB2XL U1573 ( .B0(n2055), .B1(n2183), .A0N(\register[18][24] ), .A1N(
        n2183), .Y(n650) );
  OAI2BB2XL U1574 ( .B0(n2052), .B1(n2182), .A0N(\register[18][25] ), .A1N(
        n2183), .Y(n651) );
  OAI2BB2XL U1575 ( .B0(n2049), .B1(n2182), .A0N(\register[18][26] ), .A1N(
        n2183), .Y(n652) );
  OAI2BB2XL U1576 ( .B0(n2046), .B1(n2182), .A0N(\register[18][27] ), .A1N(
        n2183), .Y(n653) );
  OAI2BB2XL U1577 ( .B0(n2043), .B1(n2181), .A0N(\register[18][28] ), .A1N(
        n2183), .Y(n654) );
  OAI2BB2XL U1578 ( .B0(n2040), .B1(n2181), .A0N(\register[18][29] ), .A1N(
        n2183), .Y(n655) );
  OAI2BB2XL U1579 ( .B0(n2037), .B1(n2181), .A0N(\register[18][30] ), .A1N(
        n2183), .Y(n656) );
  OAI2BB2XL U1580 ( .B0(n2034), .B1(n2181), .A0N(\register[18][31] ), .A1N(
        n2183), .Y(n657) );
  OAI2BB2XL U1581 ( .B0(n2127), .B1(n2177), .A0N(\register[19][0] ), .A1N(
        n2179), .Y(n658) );
  OAI2BB2XL U1582 ( .B0(n2124), .B1(n2177), .A0N(\register[19][1] ), .A1N(
        n2180), .Y(n659) );
  OAI2BB2XL U1583 ( .B0(n2121), .B1(n2177), .A0N(\register[19][2] ), .A1N(
        n2180), .Y(n660) );
  OAI2BB2XL U1584 ( .B0(n2118), .B1(n2177), .A0N(\register[19][3] ), .A1N(
        n2180), .Y(n661) );
  OAI2BB2XL U1585 ( .B0(n2115), .B1(n2177), .A0N(\register[19][4] ), .A1N(
        n2180), .Y(n662) );
  OAI2BB2XL U1586 ( .B0(n2112), .B1(n2177), .A0N(\register[19][5] ), .A1N(
        n2180), .Y(n663) );
  OAI2BB2XL U1587 ( .B0(n2109), .B1(n2177), .A0N(\register[19][6] ), .A1N(
        n2180), .Y(n664) );
  OAI2BB2XL U1588 ( .B0(n2106), .B1(n2177), .A0N(\register[19][7] ), .A1N(
        n2180), .Y(n665) );
  OAI2BB2XL U1589 ( .B0(n2103), .B1(n2178), .A0N(\register[19][8] ), .A1N(
        n2180), .Y(n666) );
  OAI2BB2XL U1590 ( .B0(n2100), .B1(n2178), .A0N(\register[19][9] ), .A1N(
        n2180), .Y(n667) );
  OAI2BB2XL U1591 ( .B0(n2097), .B1(n2178), .A0N(\register[19][10] ), .A1N(
        n2180), .Y(n668) );
  OAI2BB2XL U1592 ( .B0(n2094), .B1(n2178), .A0N(\register[19][11] ), .A1N(
        n2180), .Y(n669) );
  OAI2BB2XL U1593 ( .B0(n2091), .B1(n2178), .A0N(\register[19][12] ), .A1N(
        n2180), .Y(n670) );
  OAI2BB2XL U1594 ( .B0(n2088), .B1(n2178), .A0N(\register[19][13] ), .A1N(
        n2180), .Y(n671) );
  OAI2BB2XL U1595 ( .B0(n2085), .B1(n2178), .A0N(\register[19][14] ), .A1N(
        n2180), .Y(n672) );
  OAI2BB2XL U1596 ( .B0(n2082), .B1(n2178), .A0N(\register[19][15] ), .A1N(
        n2180), .Y(n673) );
  OAI2BB2XL U1597 ( .B0(n2079), .B1(n2179), .A0N(\register[19][16] ), .A1N(
        n2180), .Y(n674) );
  OAI2BB2XL U1598 ( .B0(n2076), .B1(n2179), .A0N(\register[19][17] ), .A1N(
        n2180), .Y(n675) );
  OAI2BB2XL U1599 ( .B0(n2073), .B1(n2178), .A0N(\register[19][18] ), .A1N(
        n2180), .Y(n676) );
  OAI2BB2XL U1600 ( .B0(n2070), .B1(n2179), .A0N(\register[19][19] ), .A1N(
        n2180), .Y(n677) );
  OAI2BB2XL U1601 ( .B0(n2067), .B1(n2179), .A0N(\register[19][20] ), .A1N(
        n2180), .Y(n678) );
  OAI2BB2XL U1602 ( .B0(n2064), .B1(n2179), .A0N(\register[19][21] ), .A1N(
        n2179), .Y(n679) );
  OAI2BB2XL U1603 ( .B0(n2061), .B1(n2179), .A0N(\register[19][22] ), .A1N(
        n2179), .Y(n680) );
  OAI2BB2XL U1604 ( .B0(n2058), .B1(n2179), .A0N(\register[19][23] ), .A1N(
        n2179), .Y(n681) );
  OAI2BB2XL U1605 ( .B0(n2055), .B1(n2179), .A0N(\register[19][24] ), .A1N(
        n2179), .Y(n682) );
  OAI2BB2XL U1606 ( .B0(n2052), .B1(n2178), .A0N(\register[19][25] ), .A1N(
        n2179), .Y(n683) );
  OAI2BB2XL U1607 ( .B0(n2049), .B1(n2178), .A0N(\register[19][26] ), .A1N(
        n2179), .Y(n684) );
  OAI2BB2XL U1608 ( .B0(n2046), .B1(n2178), .A0N(\register[19][27] ), .A1N(
        n2179), .Y(n685) );
  OAI2BB2XL U1609 ( .B0(n2043), .B1(n2177), .A0N(\register[19][28] ), .A1N(
        n2179), .Y(n686) );
  OAI2BB2XL U1610 ( .B0(n2040), .B1(n2177), .A0N(\register[19][29] ), .A1N(
        n2179), .Y(n687) );
  OAI2BB2XL U1611 ( .B0(n2037), .B1(n2177), .A0N(\register[19][30] ), .A1N(
        n2179), .Y(n688) );
  OAI2BB2XL U1612 ( .B0(n2034), .B1(n2177), .A0N(\register[19][31] ), .A1N(
        n2179), .Y(n689) );
  OAI2BB2XL U1613 ( .B0(n2126), .B1(n2173), .A0N(\register[20][0] ), .A1N(
        n2175), .Y(n690) );
  OAI2BB2XL U1614 ( .B0(n2123), .B1(n2173), .A0N(\register[20][1] ), .A1N(
        n2176), .Y(n691) );
  OAI2BB2XL U1615 ( .B0(n2120), .B1(n2173), .A0N(\register[20][2] ), .A1N(
        n2176), .Y(n692) );
  OAI2BB2XL U1616 ( .B0(n2117), .B1(n2173), .A0N(\register[20][3] ), .A1N(
        n2176), .Y(n693) );
  OAI2BB2XL U1617 ( .B0(n2114), .B1(n2173), .A0N(\register[20][4] ), .A1N(
        n2176), .Y(n694) );
  OAI2BB2XL U1618 ( .B0(n2111), .B1(n2173), .A0N(\register[20][5] ), .A1N(
        n2176), .Y(n695) );
  OAI2BB2XL U1619 ( .B0(n2108), .B1(n2173), .A0N(\register[20][6] ), .A1N(
        n2176), .Y(n696) );
  OAI2BB2XL U1620 ( .B0(n2105), .B1(n2173), .A0N(\register[20][7] ), .A1N(
        n2176), .Y(n697) );
  OAI2BB2XL U1621 ( .B0(n2102), .B1(n2174), .A0N(\register[20][8] ), .A1N(
        n2176), .Y(n698) );
  OAI2BB2XL U1622 ( .B0(n2099), .B1(n2174), .A0N(\register[20][9] ), .A1N(
        n2176), .Y(n699) );
  OAI2BB2XL U1623 ( .B0(n2096), .B1(n2174), .A0N(\register[20][10] ), .A1N(
        n2176), .Y(n700) );
  OAI2BB2XL U1624 ( .B0(n2093), .B1(n2174), .A0N(\register[20][11] ), .A1N(
        n2176), .Y(n701) );
  OAI2BB2XL U1625 ( .B0(n2090), .B1(n2174), .A0N(\register[20][12] ), .A1N(
        n2176), .Y(n702) );
  OAI2BB2XL U1626 ( .B0(n2087), .B1(n2174), .A0N(\register[20][13] ), .A1N(
        n2176), .Y(n703) );
  OAI2BB2XL U1627 ( .B0(n2084), .B1(n2174), .A0N(\register[20][14] ), .A1N(
        n2176), .Y(n704) );
  OAI2BB2XL U1628 ( .B0(n2081), .B1(n2174), .A0N(\register[20][15] ), .A1N(
        n2176), .Y(n705) );
  OAI2BB2XL U1629 ( .B0(n2078), .B1(n2175), .A0N(\register[20][16] ), .A1N(
        n2176), .Y(n706) );
  OAI2BB2XL U1630 ( .B0(n2075), .B1(n2175), .A0N(\register[20][17] ), .A1N(
        n2176), .Y(n707) );
  OAI2BB2XL U1631 ( .B0(n2072), .B1(n2174), .A0N(\register[20][18] ), .A1N(
        n2176), .Y(n708) );
  OAI2BB2XL U1632 ( .B0(n2069), .B1(n2175), .A0N(\register[20][19] ), .A1N(
        n2176), .Y(n709) );
  OAI2BB2XL U1633 ( .B0(n2066), .B1(n2175), .A0N(\register[20][20] ), .A1N(
        n2176), .Y(n710) );
  OAI2BB2XL U1634 ( .B0(n2063), .B1(n2175), .A0N(\register[20][21] ), .A1N(
        n2175), .Y(n711) );
  OAI2BB2XL U1635 ( .B0(n2060), .B1(n2175), .A0N(\register[20][22] ), .A1N(
        n2175), .Y(n712) );
  OAI2BB2XL U1636 ( .B0(n2057), .B1(n2175), .A0N(\register[20][23] ), .A1N(
        n2175), .Y(n713) );
  OAI2BB2XL U1637 ( .B0(n2054), .B1(n2175), .A0N(\register[20][24] ), .A1N(
        n2175), .Y(n714) );
  OAI2BB2XL U1638 ( .B0(n2051), .B1(n2174), .A0N(\register[20][25] ), .A1N(
        n2175), .Y(n715) );
  OAI2BB2XL U1639 ( .B0(n2048), .B1(n2174), .A0N(\register[20][26] ), .A1N(
        n2175), .Y(n716) );
  OAI2BB2XL U1640 ( .B0(n2045), .B1(n2174), .A0N(\register[20][27] ), .A1N(
        n2175), .Y(n717) );
  OAI2BB2XL U1641 ( .B0(n2042), .B1(n2173), .A0N(\register[20][28] ), .A1N(
        n2175), .Y(n718) );
  OAI2BB2XL U1642 ( .B0(n2039), .B1(n2173), .A0N(\register[20][29] ), .A1N(
        n2175), .Y(n719) );
  OAI2BB2XL U1643 ( .B0(n2036), .B1(n2173), .A0N(\register[20][30] ), .A1N(
        n2175), .Y(n720) );
  OAI2BB2XL U1644 ( .B0(n2033), .B1(n2173), .A0N(\register[20][31] ), .A1N(
        n2175), .Y(n721) );
  OAI2BB2XL U1645 ( .B0(n2126), .B1(n2169), .A0N(\register[21][0] ), .A1N(
        n2171), .Y(n722) );
  OAI2BB2XL U1646 ( .B0(n2123), .B1(n2169), .A0N(\register[21][1] ), .A1N(
        n2172), .Y(n723) );
  OAI2BB2XL U1647 ( .B0(n2120), .B1(n2169), .A0N(\register[21][2] ), .A1N(
        n2172), .Y(n724) );
  OAI2BB2XL U1648 ( .B0(n2117), .B1(n2169), .A0N(\register[21][3] ), .A1N(
        n2172), .Y(n725) );
  OAI2BB2XL U1649 ( .B0(n2114), .B1(n2169), .A0N(\register[21][4] ), .A1N(
        n2172), .Y(n726) );
  OAI2BB2XL U1650 ( .B0(n2111), .B1(n2169), .A0N(\register[21][5] ), .A1N(
        n2172), .Y(n727) );
  OAI2BB2XL U1651 ( .B0(n2108), .B1(n2169), .A0N(\register[21][6] ), .A1N(
        n2172), .Y(n728) );
  OAI2BB2XL U1652 ( .B0(n2105), .B1(n2169), .A0N(\register[21][7] ), .A1N(
        n2172), .Y(n729) );
  OAI2BB2XL U1653 ( .B0(n2102), .B1(n2170), .A0N(\register[21][8] ), .A1N(
        n2172), .Y(n730) );
  OAI2BB2XL U1654 ( .B0(n2099), .B1(n2170), .A0N(\register[21][9] ), .A1N(
        n2172), .Y(n731) );
  OAI2BB2XL U1655 ( .B0(n2096), .B1(n2170), .A0N(\register[21][10] ), .A1N(
        n2172), .Y(n732) );
  OAI2BB2XL U1656 ( .B0(n2093), .B1(n2170), .A0N(\register[21][11] ), .A1N(
        n2172), .Y(n733) );
  OAI2BB2XL U1657 ( .B0(n2090), .B1(n2170), .A0N(\register[21][12] ), .A1N(
        n2172), .Y(n734) );
  OAI2BB2XL U1658 ( .B0(n2087), .B1(n2170), .A0N(\register[21][13] ), .A1N(
        n2172), .Y(n735) );
  OAI2BB2XL U1659 ( .B0(n2084), .B1(n2170), .A0N(\register[21][14] ), .A1N(
        n2172), .Y(n736) );
  OAI2BB2XL U1660 ( .B0(n2081), .B1(n2170), .A0N(\register[21][15] ), .A1N(
        n2172), .Y(n737) );
  OAI2BB2XL U1661 ( .B0(n2078), .B1(n2171), .A0N(\register[21][16] ), .A1N(
        n2172), .Y(n738) );
  OAI2BB2XL U1662 ( .B0(n2075), .B1(n2171), .A0N(\register[21][17] ), .A1N(
        n2172), .Y(n739) );
  OAI2BB2XL U1663 ( .B0(n2072), .B1(n2170), .A0N(\register[21][18] ), .A1N(
        n2172), .Y(n740) );
  OAI2BB2XL U1664 ( .B0(n2069), .B1(n2171), .A0N(\register[21][19] ), .A1N(
        n2172), .Y(n741) );
  OAI2BB2XL U1665 ( .B0(n2066), .B1(n2171), .A0N(\register[21][20] ), .A1N(
        n2172), .Y(n742) );
  OAI2BB2XL U1666 ( .B0(n2063), .B1(n2171), .A0N(\register[21][21] ), .A1N(
        n2171), .Y(n743) );
  OAI2BB2XL U1667 ( .B0(n2060), .B1(n2171), .A0N(\register[21][22] ), .A1N(
        n2171), .Y(n744) );
  OAI2BB2XL U1668 ( .B0(n2057), .B1(n2171), .A0N(\register[21][23] ), .A1N(
        n2171), .Y(n745) );
  OAI2BB2XL U1669 ( .B0(n2054), .B1(n2171), .A0N(\register[21][24] ), .A1N(
        n2171), .Y(n746) );
  OAI2BB2XL U1670 ( .B0(n2051), .B1(n2170), .A0N(\register[21][25] ), .A1N(
        n2171), .Y(n747) );
  OAI2BB2XL U1671 ( .B0(n2048), .B1(n2170), .A0N(\register[21][26] ), .A1N(
        n2171), .Y(n748) );
  OAI2BB2XL U1672 ( .B0(n2045), .B1(n2170), .A0N(\register[21][27] ), .A1N(
        n2171), .Y(n749) );
  OAI2BB2XL U1673 ( .B0(n2042), .B1(n2169), .A0N(\register[21][28] ), .A1N(
        n2171), .Y(n750) );
  OAI2BB2XL U1674 ( .B0(n2039), .B1(n2169), .A0N(\register[21][29] ), .A1N(
        n2171), .Y(n751) );
  OAI2BB2XL U1675 ( .B0(n2036), .B1(n2169), .A0N(\register[21][30] ), .A1N(
        n2171), .Y(n752) );
  OAI2BB2XL U1676 ( .B0(n2033), .B1(n2169), .A0N(\register[21][31] ), .A1N(
        n2171), .Y(n753) );
  OAI2BB2XL U1677 ( .B0(n2126), .B1(n2165), .A0N(\register[22][0] ), .A1N(
        n2167), .Y(n754) );
  OAI2BB2XL U1678 ( .B0(n2123), .B1(n2165), .A0N(\register[22][1] ), .A1N(
        n2168), .Y(n755) );
  OAI2BB2XL U1679 ( .B0(n2120), .B1(n2165), .A0N(\register[22][2] ), .A1N(
        n2168), .Y(n756) );
  OAI2BB2XL U1680 ( .B0(n2117), .B1(n2165), .A0N(\register[22][3] ), .A1N(
        n2168), .Y(n757) );
  OAI2BB2XL U1681 ( .B0(n2114), .B1(n2165), .A0N(\register[22][4] ), .A1N(
        n2168), .Y(n758) );
  OAI2BB2XL U1682 ( .B0(n2111), .B1(n2165), .A0N(\register[22][5] ), .A1N(
        n2168), .Y(n759) );
  OAI2BB2XL U1683 ( .B0(n2108), .B1(n2165), .A0N(\register[22][6] ), .A1N(
        n2168), .Y(n760) );
  OAI2BB2XL U1684 ( .B0(n2105), .B1(n2165), .A0N(\register[22][7] ), .A1N(
        n2168), .Y(n761) );
  OAI2BB2XL U1685 ( .B0(n2102), .B1(n2166), .A0N(\register[22][8] ), .A1N(
        n2168), .Y(n762) );
  OAI2BB2XL U1686 ( .B0(n2099), .B1(n2166), .A0N(\register[22][9] ), .A1N(
        n2168), .Y(n763) );
  OAI2BB2XL U1687 ( .B0(n2096), .B1(n2166), .A0N(\register[22][10] ), .A1N(
        n2168), .Y(n764) );
  OAI2BB2XL U1688 ( .B0(n2093), .B1(n2166), .A0N(\register[22][11] ), .A1N(
        n2168), .Y(n765) );
  OAI2BB2XL U1689 ( .B0(n2090), .B1(n2166), .A0N(\register[22][12] ), .A1N(
        n2168), .Y(n766) );
  OAI2BB2XL U1690 ( .B0(n2087), .B1(n2166), .A0N(\register[22][13] ), .A1N(
        n2168), .Y(n767) );
  OAI2BB2XL U1691 ( .B0(n2084), .B1(n2166), .A0N(\register[22][14] ), .A1N(
        n2168), .Y(n768) );
  OAI2BB2XL U1692 ( .B0(n2081), .B1(n2166), .A0N(\register[22][15] ), .A1N(
        n2168), .Y(n769) );
  OAI2BB2XL U1693 ( .B0(n2078), .B1(n2167), .A0N(\register[22][16] ), .A1N(
        n2168), .Y(n770) );
  OAI2BB2XL U1694 ( .B0(n2075), .B1(n2167), .A0N(\register[22][17] ), .A1N(
        n2168), .Y(n771) );
  OAI2BB2XL U1695 ( .B0(n2072), .B1(n2166), .A0N(\register[22][18] ), .A1N(
        n2168), .Y(n772) );
  OAI2BB2XL U1696 ( .B0(n2069), .B1(n2167), .A0N(\register[22][19] ), .A1N(
        n2168), .Y(n773) );
  OAI2BB2XL U1697 ( .B0(n2066), .B1(n2167), .A0N(\register[22][20] ), .A1N(
        n2168), .Y(n774) );
  OAI2BB2XL U1698 ( .B0(n2063), .B1(n2167), .A0N(\register[22][21] ), .A1N(
        n2167), .Y(n775) );
  OAI2BB2XL U1699 ( .B0(n2060), .B1(n2167), .A0N(\register[22][22] ), .A1N(
        n2167), .Y(n776) );
  OAI2BB2XL U1700 ( .B0(n2057), .B1(n2167), .A0N(\register[22][23] ), .A1N(
        n2167), .Y(n777) );
  OAI2BB2XL U1701 ( .B0(n2054), .B1(n2167), .A0N(\register[22][24] ), .A1N(
        n2167), .Y(n778) );
  OAI2BB2XL U1702 ( .B0(n2051), .B1(n2166), .A0N(\register[22][25] ), .A1N(
        n2167), .Y(n779) );
  OAI2BB2XL U1703 ( .B0(n2048), .B1(n2166), .A0N(\register[22][26] ), .A1N(
        n2167), .Y(n780) );
  OAI2BB2XL U1704 ( .B0(n2045), .B1(n2166), .A0N(\register[22][27] ), .A1N(
        n2167), .Y(n781) );
  OAI2BB2XL U1705 ( .B0(n2042), .B1(n2165), .A0N(\register[22][28] ), .A1N(
        n2167), .Y(n782) );
  OAI2BB2XL U1706 ( .B0(n2039), .B1(n2165), .A0N(\register[22][29] ), .A1N(
        n2167), .Y(n783) );
  OAI2BB2XL U1707 ( .B0(n2036), .B1(n2165), .A0N(\register[22][30] ), .A1N(
        n2167), .Y(n784) );
  OAI2BB2XL U1708 ( .B0(n2033), .B1(n2165), .A0N(\register[22][31] ), .A1N(
        n2167), .Y(n785) );
  OAI2BB2XL U1709 ( .B0(n2126), .B1(n2161), .A0N(\register[23][0] ), .A1N(
        n2163), .Y(n786) );
  OAI2BB2XL U1710 ( .B0(n2123), .B1(n2161), .A0N(\register[23][1] ), .A1N(
        n2164), .Y(n787) );
  OAI2BB2XL U1711 ( .B0(n2120), .B1(n2161), .A0N(\register[23][2] ), .A1N(
        n2164), .Y(n788) );
  OAI2BB2XL U1712 ( .B0(n2117), .B1(n2161), .A0N(\register[23][3] ), .A1N(
        n2164), .Y(n789) );
  OAI2BB2XL U1713 ( .B0(n2114), .B1(n2161), .A0N(\register[23][4] ), .A1N(
        n2164), .Y(n790) );
  OAI2BB2XL U1714 ( .B0(n2111), .B1(n2161), .A0N(\register[23][5] ), .A1N(
        n2164), .Y(n791) );
  OAI2BB2XL U1715 ( .B0(n2108), .B1(n2161), .A0N(\register[23][6] ), .A1N(
        n2164), .Y(n792) );
  OAI2BB2XL U1716 ( .B0(n2105), .B1(n2161), .A0N(\register[23][7] ), .A1N(
        n2164), .Y(n793) );
  OAI2BB2XL U1717 ( .B0(n2102), .B1(n2162), .A0N(\register[23][8] ), .A1N(
        n2164), .Y(n794) );
  OAI2BB2XL U1718 ( .B0(n2099), .B1(n2162), .A0N(\register[23][9] ), .A1N(
        n2164), .Y(n795) );
  OAI2BB2XL U1719 ( .B0(n2096), .B1(n2162), .A0N(\register[23][10] ), .A1N(
        n2164), .Y(n796) );
  OAI2BB2XL U1720 ( .B0(n2093), .B1(n2162), .A0N(\register[23][11] ), .A1N(
        n2164), .Y(n797) );
  OAI2BB2XL U1721 ( .B0(n2090), .B1(n2162), .A0N(\register[23][12] ), .A1N(
        n2164), .Y(n798) );
  OAI2BB2XL U1722 ( .B0(n2087), .B1(n2162), .A0N(\register[23][13] ), .A1N(
        n2164), .Y(n799) );
  OAI2BB2XL U1723 ( .B0(n2084), .B1(n2162), .A0N(\register[23][14] ), .A1N(
        n2164), .Y(n800) );
  OAI2BB2XL U1724 ( .B0(n2081), .B1(n2162), .A0N(\register[23][15] ), .A1N(
        n2164), .Y(n801) );
  OAI2BB2XL U1725 ( .B0(n2078), .B1(n2163), .A0N(\register[23][16] ), .A1N(
        n2164), .Y(n802) );
  OAI2BB2XL U1726 ( .B0(n2075), .B1(n2163), .A0N(\register[23][17] ), .A1N(
        n2164), .Y(n803) );
  OAI2BB2XL U1727 ( .B0(n2072), .B1(n2162), .A0N(\register[23][18] ), .A1N(
        n2164), .Y(n804) );
  OAI2BB2XL U1728 ( .B0(n2069), .B1(n2163), .A0N(\register[23][19] ), .A1N(
        n2164), .Y(n805) );
  OAI2BB2XL U1729 ( .B0(n2066), .B1(n2163), .A0N(\register[23][20] ), .A1N(
        n2164), .Y(n806) );
  OAI2BB2XL U1730 ( .B0(n2063), .B1(n2163), .A0N(\register[23][21] ), .A1N(
        n2163), .Y(n807) );
  OAI2BB2XL U1731 ( .B0(n2060), .B1(n2163), .A0N(\register[23][22] ), .A1N(
        n2163), .Y(n808) );
  OAI2BB2XL U1732 ( .B0(n2057), .B1(n2163), .A0N(\register[23][23] ), .A1N(
        n2163), .Y(n809) );
  OAI2BB2XL U1733 ( .B0(n2054), .B1(n2163), .A0N(\register[23][24] ), .A1N(
        n2163), .Y(n810) );
  OAI2BB2XL U1734 ( .B0(n2051), .B1(n2162), .A0N(\register[23][25] ), .A1N(
        n2163), .Y(n811) );
  OAI2BB2XL U1735 ( .B0(n2048), .B1(n2162), .A0N(\register[23][26] ), .A1N(
        n2163), .Y(n812) );
  OAI2BB2XL U1736 ( .B0(n2045), .B1(n2162), .A0N(\register[23][27] ), .A1N(
        n2163), .Y(n813) );
  OAI2BB2XL U1737 ( .B0(n2042), .B1(n2161), .A0N(\register[23][28] ), .A1N(
        n2163), .Y(n814) );
  OAI2BB2XL U1738 ( .B0(n2039), .B1(n2161), .A0N(\register[23][29] ), .A1N(
        n2163), .Y(n815) );
  OAI2BB2XL U1739 ( .B0(n2036), .B1(n2161), .A0N(\register[23][30] ), .A1N(
        n2163), .Y(n816) );
  OAI2BB2XL U1740 ( .B0(n2033), .B1(n2161), .A0N(\register[23][31] ), .A1N(
        n2163), .Y(n817) );
  OAI2BB2XL U1741 ( .B0(n2126), .B1(n2157), .A0N(\register[24][0] ), .A1N(
        n2159), .Y(n818) );
  OAI2BB2XL U1742 ( .B0(n2123), .B1(n2157), .A0N(\register[24][1] ), .A1N(
        n2160), .Y(n819) );
  OAI2BB2XL U1743 ( .B0(n2120), .B1(n2157), .A0N(\register[24][2] ), .A1N(
        n2160), .Y(n820) );
  OAI2BB2XL U1744 ( .B0(n2117), .B1(n2157), .A0N(\register[24][3] ), .A1N(
        n2160), .Y(n821) );
  OAI2BB2XL U1745 ( .B0(n2114), .B1(n2157), .A0N(\register[24][4] ), .A1N(
        n2160), .Y(n822) );
  OAI2BB2XL U1746 ( .B0(n2111), .B1(n2157), .A0N(\register[24][5] ), .A1N(
        n2160), .Y(n823) );
  OAI2BB2XL U1747 ( .B0(n2108), .B1(n2157), .A0N(\register[24][6] ), .A1N(
        n2160), .Y(n824) );
  OAI2BB2XL U1748 ( .B0(n2105), .B1(n2157), .A0N(\register[24][7] ), .A1N(
        n2160), .Y(n825) );
  OAI2BB2XL U1749 ( .B0(n2102), .B1(n2158), .A0N(\register[24][8] ), .A1N(
        n2160), .Y(n826) );
  OAI2BB2XL U1750 ( .B0(n2099), .B1(n2158), .A0N(\register[24][9] ), .A1N(
        n2160), .Y(n827) );
  OAI2BB2XL U1751 ( .B0(n2096), .B1(n2158), .A0N(\register[24][10] ), .A1N(
        n2160), .Y(n828) );
  OAI2BB2XL U1752 ( .B0(n2093), .B1(n2158), .A0N(\register[24][11] ), .A1N(
        n2160), .Y(n829) );
  OAI2BB2XL U1753 ( .B0(n2090), .B1(n2158), .A0N(\register[24][12] ), .A1N(
        n2160), .Y(n830) );
  OAI2BB2XL U1754 ( .B0(n2087), .B1(n2158), .A0N(\register[24][13] ), .A1N(
        n2160), .Y(n831) );
  OAI2BB2XL U1755 ( .B0(n2084), .B1(n2158), .A0N(\register[24][14] ), .A1N(
        n2160), .Y(n832) );
  OAI2BB2XL U1756 ( .B0(n2081), .B1(n2158), .A0N(\register[24][15] ), .A1N(
        n2160), .Y(n833) );
  OAI2BB2XL U1757 ( .B0(n2078), .B1(n2159), .A0N(\register[24][16] ), .A1N(
        n2160), .Y(n834) );
  OAI2BB2XL U1758 ( .B0(n2075), .B1(n2159), .A0N(\register[24][17] ), .A1N(
        n2160), .Y(n835) );
  OAI2BB2XL U1759 ( .B0(n2072), .B1(n2158), .A0N(\register[24][18] ), .A1N(
        n2160), .Y(n836) );
  OAI2BB2XL U1760 ( .B0(n2069), .B1(n2159), .A0N(\register[24][19] ), .A1N(
        n2160), .Y(n837) );
  OAI2BB2XL U1761 ( .B0(n2066), .B1(n2159), .A0N(\register[24][20] ), .A1N(
        n2160), .Y(n838) );
  OAI2BB2XL U1762 ( .B0(n2063), .B1(n2159), .A0N(\register[24][21] ), .A1N(
        n2159), .Y(n839) );
  OAI2BB2XL U1763 ( .B0(n2060), .B1(n2159), .A0N(\register[24][22] ), .A1N(
        n2159), .Y(n840) );
  OAI2BB2XL U1764 ( .B0(n2057), .B1(n2159), .A0N(\register[24][23] ), .A1N(
        n2159), .Y(n841) );
  OAI2BB2XL U1765 ( .B0(n2054), .B1(n2159), .A0N(\register[24][24] ), .A1N(
        n2159), .Y(n842) );
  OAI2BB2XL U1766 ( .B0(n2051), .B1(n2158), .A0N(\register[24][25] ), .A1N(
        n2159), .Y(n843) );
  OAI2BB2XL U1767 ( .B0(n2048), .B1(n2158), .A0N(\register[24][26] ), .A1N(
        n2159), .Y(n844) );
  OAI2BB2XL U1768 ( .B0(n2045), .B1(n2158), .A0N(\register[24][27] ), .A1N(
        n2159), .Y(n845) );
  OAI2BB2XL U1769 ( .B0(n2042), .B1(n2157), .A0N(\register[24][28] ), .A1N(
        n2159), .Y(n846) );
  OAI2BB2XL U1770 ( .B0(n2039), .B1(n2157), .A0N(\register[24][29] ), .A1N(
        n2159), .Y(n847) );
  OAI2BB2XL U1771 ( .B0(n2036), .B1(n2157), .A0N(\register[24][30] ), .A1N(
        n2159), .Y(n848) );
  OAI2BB2XL U1772 ( .B0(n2033), .B1(n2157), .A0N(\register[24][31] ), .A1N(
        n2159), .Y(n849) );
  OAI2BB2XL U1773 ( .B0(n2126), .B1(n2153), .A0N(\register[25][0] ), .A1N(
        n2155), .Y(n850) );
  OAI2BB2XL U1774 ( .B0(n2123), .B1(n2153), .A0N(\register[25][1] ), .A1N(
        n2156), .Y(n851) );
  OAI2BB2XL U1775 ( .B0(n2120), .B1(n2153), .A0N(\register[25][2] ), .A1N(
        n2156), .Y(n852) );
  OAI2BB2XL U1776 ( .B0(n2117), .B1(n2153), .A0N(\register[25][3] ), .A1N(
        n2156), .Y(n853) );
  OAI2BB2XL U1777 ( .B0(n2114), .B1(n2153), .A0N(\register[25][4] ), .A1N(
        n2156), .Y(n854) );
  OAI2BB2XL U1778 ( .B0(n2111), .B1(n2153), .A0N(\register[25][5] ), .A1N(
        n2156), .Y(n855) );
  OAI2BB2XL U1779 ( .B0(n2108), .B1(n2153), .A0N(\register[25][6] ), .A1N(
        n2156), .Y(n856) );
  OAI2BB2XL U1780 ( .B0(n2105), .B1(n2153), .A0N(\register[25][7] ), .A1N(
        n2156), .Y(n857) );
  OAI2BB2XL U1781 ( .B0(n2102), .B1(n2154), .A0N(\register[25][8] ), .A1N(
        n2156), .Y(n858) );
  OAI2BB2XL U1782 ( .B0(n2099), .B1(n2154), .A0N(\register[25][9] ), .A1N(
        n2156), .Y(n859) );
  OAI2BB2XL U1783 ( .B0(n2096), .B1(n2154), .A0N(\register[25][10] ), .A1N(
        n2156), .Y(n860) );
  OAI2BB2XL U1784 ( .B0(n2093), .B1(n2154), .A0N(\register[25][11] ), .A1N(
        n2156), .Y(n861) );
  OAI2BB2XL U1785 ( .B0(n2090), .B1(n2154), .A0N(\register[25][12] ), .A1N(
        n2156), .Y(n862) );
  OAI2BB2XL U1786 ( .B0(n2087), .B1(n2154), .A0N(\register[25][13] ), .A1N(
        n2156), .Y(n863) );
  OAI2BB2XL U1787 ( .B0(n2084), .B1(n2154), .A0N(\register[25][14] ), .A1N(
        n2156), .Y(n864) );
  OAI2BB2XL U1788 ( .B0(n2081), .B1(n2154), .A0N(\register[25][15] ), .A1N(
        n2156), .Y(n865) );
  OAI2BB2XL U1789 ( .B0(n2078), .B1(n2155), .A0N(\register[25][16] ), .A1N(
        n2156), .Y(n866) );
  OAI2BB2XL U1790 ( .B0(n2075), .B1(n2155), .A0N(\register[25][17] ), .A1N(
        n2156), .Y(n867) );
  OAI2BB2XL U1791 ( .B0(n2072), .B1(n2154), .A0N(\register[25][18] ), .A1N(
        n2156), .Y(n868) );
  OAI2BB2XL U1792 ( .B0(n2069), .B1(n2155), .A0N(\register[25][19] ), .A1N(
        n2156), .Y(n869) );
  OAI2BB2XL U1793 ( .B0(n2066), .B1(n2155), .A0N(\register[25][20] ), .A1N(
        n2156), .Y(n870) );
  OAI2BB2XL U1794 ( .B0(n2063), .B1(n2155), .A0N(\register[25][21] ), .A1N(
        n2155), .Y(n871) );
  OAI2BB2XL U1795 ( .B0(n2060), .B1(n2155), .A0N(\register[25][22] ), .A1N(
        n2155), .Y(n872) );
  OAI2BB2XL U1796 ( .B0(n2057), .B1(n2155), .A0N(\register[25][23] ), .A1N(
        n2155), .Y(n873) );
  OAI2BB2XL U1797 ( .B0(n2054), .B1(n2155), .A0N(\register[25][24] ), .A1N(
        n2155), .Y(n874) );
  OAI2BB2XL U1798 ( .B0(n2051), .B1(n2154), .A0N(\register[25][25] ), .A1N(
        n2155), .Y(n875) );
  OAI2BB2XL U1799 ( .B0(n2048), .B1(n2154), .A0N(\register[25][26] ), .A1N(
        n2155), .Y(n876) );
  OAI2BB2XL U1800 ( .B0(n2045), .B1(n2154), .A0N(\register[25][27] ), .A1N(
        n2155), .Y(n877) );
  OAI2BB2XL U1801 ( .B0(n2042), .B1(n2153), .A0N(\register[25][28] ), .A1N(
        n2155), .Y(n878) );
  OAI2BB2XL U1802 ( .B0(n2039), .B1(n2153), .A0N(\register[25][29] ), .A1N(
        n2155), .Y(n879) );
  OAI2BB2XL U1803 ( .B0(n2036), .B1(n2153), .A0N(\register[25][30] ), .A1N(
        n2155), .Y(n880) );
  OAI2BB2XL U1804 ( .B0(n2033), .B1(n2153), .A0N(\register[25][31] ), .A1N(
        n2155), .Y(n881) );
  OAI2BB2XL U1805 ( .B0(n2126), .B1(n2149), .A0N(\register[26][0] ), .A1N(
        n2151), .Y(n882) );
  OAI2BB2XL U1806 ( .B0(n2123), .B1(n2149), .A0N(\register[26][1] ), .A1N(
        n2152), .Y(n883) );
  OAI2BB2XL U1807 ( .B0(n2120), .B1(n2149), .A0N(\register[26][2] ), .A1N(
        n2152), .Y(n884) );
  OAI2BB2XL U1808 ( .B0(n2117), .B1(n2149), .A0N(\register[26][3] ), .A1N(
        n2152), .Y(n885) );
  OAI2BB2XL U1809 ( .B0(n2114), .B1(n2149), .A0N(\register[26][4] ), .A1N(
        n2152), .Y(n886) );
  OAI2BB2XL U1810 ( .B0(n2111), .B1(n2149), .A0N(\register[26][5] ), .A1N(
        n2152), .Y(n887) );
  OAI2BB2XL U1811 ( .B0(n2108), .B1(n2149), .A0N(\register[26][6] ), .A1N(
        n2152), .Y(n888) );
  OAI2BB2XL U1812 ( .B0(n2105), .B1(n2149), .A0N(\register[26][7] ), .A1N(
        n2152), .Y(n889) );
  OAI2BB2XL U1813 ( .B0(n2102), .B1(n2150), .A0N(\register[26][8] ), .A1N(
        n2152), .Y(n890) );
  OAI2BB2XL U1814 ( .B0(n2099), .B1(n2150), .A0N(\register[26][9] ), .A1N(
        n2152), .Y(n891) );
  OAI2BB2XL U1815 ( .B0(n2096), .B1(n2150), .A0N(\register[26][10] ), .A1N(
        n2152), .Y(n892) );
  OAI2BB2XL U1816 ( .B0(n2093), .B1(n2150), .A0N(\register[26][11] ), .A1N(
        n2152), .Y(n893) );
  OAI2BB2XL U1817 ( .B0(n2090), .B1(n2150), .A0N(\register[26][12] ), .A1N(
        n2152), .Y(n894) );
  OAI2BB2XL U1818 ( .B0(n2087), .B1(n2150), .A0N(\register[26][13] ), .A1N(
        n2152), .Y(n895) );
  OAI2BB2XL U1819 ( .B0(n2084), .B1(n2150), .A0N(\register[26][14] ), .A1N(
        n2152), .Y(n896) );
  OAI2BB2XL U1820 ( .B0(n2081), .B1(n2150), .A0N(\register[26][15] ), .A1N(
        n2152), .Y(n897) );
  OAI2BB2XL U1821 ( .B0(n2078), .B1(n2151), .A0N(\register[26][16] ), .A1N(
        n2152), .Y(n898) );
  OAI2BB2XL U1822 ( .B0(n2075), .B1(n2151), .A0N(\register[26][17] ), .A1N(
        n2152), .Y(n899) );
  OAI2BB2XL U1823 ( .B0(n2072), .B1(n2150), .A0N(\register[26][18] ), .A1N(
        n2152), .Y(n900) );
  OAI2BB2XL U1824 ( .B0(n2069), .B1(n2151), .A0N(\register[26][19] ), .A1N(
        n2152), .Y(n901) );
  OAI2BB2XL U1825 ( .B0(n2066), .B1(n2151), .A0N(\register[26][20] ), .A1N(
        n2152), .Y(n902) );
  OAI2BB2XL U1826 ( .B0(n2063), .B1(n2151), .A0N(\register[26][21] ), .A1N(
        n2151), .Y(n903) );
  OAI2BB2XL U1827 ( .B0(n2060), .B1(n2151), .A0N(\register[26][22] ), .A1N(
        n2151), .Y(n904) );
  OAI2BB2XL U1828 ( .B0(n2057), .B1(n2151), .A0N(\register[26][23] ), .A1N(
        n2151), .Y(n905) );
  OAI2BB2XL U1829 ( .B0(n2054), .B1(n2151), .A0N(\register[26][24] ), .A1N(
        n2151), .Y(n906) );
  OAI2BB2XL U1830 ( .B0(n2051), .B1(n2150), .A0N(\register[26][25] ), .A1N(
        n2151), .Y(n907) );
  OAI2BB2XL U1831 ( .B0(n2048), .B1(n2150), .A0N(\register[26][26] ), .A1N(
        n2151), .Y(n908) );
  OAI2BB2XL U1832 ( .B0(n2045), .B1(n2150), .A0N(\register[26][27] ), .A1N(
        n2151), .Y(n909) );
  OAI2BB2XL U1833 ( .B0(n2042), .B1(n2149), .A0N(\register[26][28] ), .A1N(
        n2151), .Y(n910) );
  OAI2BB2XL U1834 ( .B0(n2039), .B1(n2149), .A0N(\register[26][29] ), .A1N(
        n2151), .Y(n911) );
  OAI2BB2XL U1835 ( .B0(n2036), .B1(n2149), .A0N(\register[26][30] ), .A1N(
        n2151), .Y(n912) );
  OAI2BB2XL U1836 ( .B0(n2033), .B1(n2149), .A0N(\register[26][31] ), .A1N(
        n2151), .Y(n913) );
  OAI2BB2XL U1837 ( .B0(n2126), .B1(n2145), .A0N(\register[27][0] ), .A1N(
        n2147), .Y(n914) );
  OAI2BB2XL U1838 ( .B0(n2123), .B1(n2145), .A0N(\register[27][1] ), .A1N(
        n2148), .Y(n915) );
  OAI2BB2XL U1839 ( .B0(n2120), .B1(n2145), .A0N(\register[27][2] ), .A1N(
        n2148), .Y(n916) );
  OAI2BB2XL U1840 ( .B0(n2117), .B1(n2145), .A0N(\register[27][3] ), .A1N(
        n2148), .Y(n917) );
  OAI2BB2XL U1841 ( .B0(n2114), .B1(n2145), .A0N(\register[27][4] ), .A1N(
        n2148), .Y(n918) );
  OAI2BB2XL U1842 ( .B0(n2111), .B1(n2145), .A0N(\register[27][5] ), .A1N(
        n2148), .Y(n919) );
  OAI2BB2XL U1843 ( .B0(n2108), .B1(n2145), .A0N(\register[27][6] ), .A1N(
        n2148), .Y(n920) );
  OAI2BB2XL U1844 ( .B0(n2105), .B1(n2145), .A0N(\register[27][7] ), .A1N(
        n2148), .Y(n921) );
  OAI2BB2XL U1845 ( .B0(n2102), .B1(n2146), .A0N(\register[27][8] ), .A1N(
        n2148), .Y(n922) );
  OAI2BB2XL U1846 ( .B0(n2099), .B1(n2146), .A0N(\register[27][9] ), .A1N(
        n2148), .Y(n923) );
  OAI2BB2XL U1847 ( .B0(n2096), .B1(n2146), .A0N(\register[27][10] ), .A1N(
        n2148), .Y(n924) );
  OAI2BB2XL U1848 ( .B0(n2093), .B1(n2146), .A0N(\register[27][11] ), .A1N(
        n2148), .Y(n925) );
  OAI2BB2XL U1849 ( .B0(n2090), .B1(n2146), .A0N(\register[27][12] ), .A1N(
        n2148), .Y(n926) );
  OAI2BB2XL U1850 ( .B0(n2087), .B1(n2146), .A0N(\register[27][13] ), .A1N(
        n2148), .Y(n927) );
  OAI2BB2XL U1851 ( .B0(n2084), .B1(n2146), .A0N(\register[27][14] ), .A1N(
        n2148), .Y(n928) );
  OAI2BB2XL U1852 ( .B0(n2081), .B1(n2146), .A0N(\register[27][15] ), .A1N(
        n2148), .Y(n929) );
  OAI2BB2XL U1853 ( .B0(n2078), .B1(n2147), .A0N(\register[27][16] ), .A1N(
        n2148), .Y(n930) );
  OAI2BB2XL U1854 ( .B0(n2075), .B1(n2147), .A0N(\register[27][17] ), .A1N(
        n2148), .Y(n931) );
  OAI2BB2XL U1855 ( .B0(n2072), .B1(n2146), .A0N(\register[27][18] ), .A1N(
        n2148), .Y(n932) );
  OAI2BB2XL U1856 ( .B0(n2069), .B1(n2147), .A0N(\register[27][19] ), .A1N(
        n2148), .Y(n933) );
  OAI2BB2XL U1857 ( .B0(n2066), .B1(n2147), .A0N(\register[27][20] ), .A1N(
        n2148), .Y(n934) );
  OAI2BB2XL U1858 ( .B0(n2063), .B1(n2147), .A0N(\register[27][21] ), .A1N(
        n2147), .Y(n935) );
  OAI2BB2XL U1859 ( .B0(n2060), .B1(n2147), .A0N(\register[27][22] ), .A1N(
        n2147), .Y(n936) );
  OAI2BB2XL U1860 ( .B0(n2057), .B1(n2147), .A0N(\register[27][23] ), .A1N(
        n2147), .Y(n937) );
  OAI2BB2XL U1861 ( .B0(n2054), .B1(n2147), .A0N(\register[27][24] ), .A1N(
        n2147), .Y(n938) );
  OAI2BB2XL U1862 ( .B0(n2051), .B1(n2146), .A0N(\register[27][25] ), .A1N(
        n2147), .Y(n939) );
  OAI2BB2XL U1863 ( .B0(n2048), .B1(n2146), .A0N(\register[27][26] ), .A1N(
        n2147), .Y(n940) );
  OAI2BB2XL U1864 ( .B0(n2045), .B1(n2146), .A0N(\register[27][27] ), .A1N(
        n2147), .Y(n941) );
  OAI2BB2XL U1865 ( .B0(n2042), .B1(n2145), .A0N(\register[27][28] ), .A1N(
        n2147), .Y(n942) );
  OAI2BB2XL U1866 ( .B0(n2039), .B1(n2145), .A0N(\register[27][29] ), .A1N(
        n2147), .Y(n943) );
  OAI2BB2XL U1867 ( .B0(n2036), .B1(n2145), .A0N(\register[27][30] ), .A1N(
        n2147), .Y(n944) );
  OAI2BB2XL U1868 ( .B0(n2033), .B1(n2145), .A0N(\register[27][31] ), .A1N(
        n2147), .Y(n945) );
  OAI2BB2XL U1869 ( .B0(n2126), .B1(n2141), .A0N(\register[28][0] ), .A1N(
        n2143), .Y(n946) );
  OAI2BB2XL U1870 ( .B0(n2123), .B1(n2141), .A0N(\register[28][1] ), .A1N(
        n2144), .Y(n947) );
  OAI2BB2XL U1871 ( .B0(n2120), .B1(n2141), .A0N(\register[28][2] ), .A1N(
        n2144), .Y(n948) );
  OAI2BB2XL U1872 ( .B0(n2117), .B1(n2141), .A0N(\register[28][3] ), .A1N(
        n2144), .Y(n949) );
  OAI2BB2XL U1873 ( .B0(n2114), .B1(n2141), .A0N(\register[28][4] ), .A1N(
        n2144), .Y(n950) );
  OAI2BB2XL U1874 ( .B0(n2111), .B1(n2141), .A0N(\register[28][5] ), .A1N(
        n2144), .Y(n951) );
  OAI2BB2XL U1875 ( .B0(n2108), .B1(n2141), .A0N(\register[28][6] ), .A1N(
        n2144), .Y(n952) );
  OAI2BB2XL U1876 ( .B0(n2105), .B1(n2141), .A0N(\register[28][7] ), .A1N(
        n2144), .Y(n953) );
  OAI2BB2XL U1877 ( .B0(n2102), .B1(n2142), .A0N(\register[28][8] ), .A1N(
        n2144), .Y(n954) );
  OAI2BB2XL U1878 ( .B0(n2099), .B1(n2142), .A0N(\register[28][9] ), .A1N(
        n2144), .Y(n955) );
  OAI2BB2XL U1879 ( .B0(n2096), .B1(n2142), .A0N(\register[28][10] ), .A1N(
        n2144), .Y(n956) );
  OAI2BB2XL U1880 ( .B0(n2093), .B1(n2142), .A0N(\register[28][11] ), .A1N(
        n2144), .Y(n957) );
  OAI2BB2XL U1881 ( .B0(n2090), .B1(n2142), .A0N(\register[28][12] ), .A1N(
        n2144), .Y(n958) );
  OAI2BB2XL U1882 ( .B0(n2087), .B1(n2142), .A0N(\register[28][13] ), .A1N(
        n2144), .Y(n959) );
  OAI2BB2XL U1883 ( .B0(n2084), .B1(n2142), .A0N(\register[28][14] ), .A1N(
        n2144), .Y(n960) );
  OAI2BB2XL U1884 ( .B0(n2081), .B1(n2142), .A0N(\register[28][15] ), .A1N(
        n2144), .Y(n961) );
  OAI2BB2XL U1885 ( .B0(n2078), .B1(n2143), .A0N(\register[28][16] ), .A1N(
        n2144), .Y(n962) );
  OAI2BB2XL U1886 ( .B0(n2075), .B1(n2143), .A0N(\register[28][17] ), .A1N(
        n2144), .Y(n963) );
  OAI2BB2XL U1887 ( .B0(n2072), .B1(n2142), .A0N(\register[28][18] ), .A1N(
        n2144), .Y(n964) );
  OAI2BB2XL U1888 ( .B0(n2069), .B1(n2143), .A0N(\register[28][19] ), .A1N(
        n2144), .Y(n965) );
  OAI2BB2XL U1889 ( .B0(n2066), .B1(n2143), .A0N(\register[28][20] ), .A1N(
        n2144), .Y(n966) );
  OAI2BB2XL U1890 ( .B0(n2063), .B1(n2143), .A0N(\register[28][21] ), .A1N(
        n2143), .Y(n967) );
  OAI2BB2XL U1891 ( .B0(n2060), .B1(n2143), .A0N(\register[28][22] ), .A1N(
        n2143), .Y(n968) );
  OAI2BB2XL U1892 ( .B0(n2057), .B1(n2143), .A0N(\register[28][23] ), .A1N(
        n2143), .Y(n969) );
  OAI2BB2XL U1893 ( .B0(n2054), .B1(n2143), .A0N(\register[28][24] ), .A1N(
        n2143), .Y(n970) );
  OAI2BB2XL U1894 ( .B0(n2051), .B1(n2142), .A0N(\register[28][25] ), .A1N(
        n2143), .Y(n971) );
  OAI2BB2XL U1895 ( .B0(n2048), .B1(n2142), .A0N(\register[28][26] ), .A1N(
        n2143), .Y(n972) );
  OAI2BB2XL U1896 ( .B0(n2045), .B1(n2142), .A0N(\register[28][27] ), .A1N(
        n2143), .Y(n973) );
  OAI2BB2XL U1897 ( .B0(n2042), .B1(n2141), .A0N(\register[28][28] ), .A1N(
        n2143), .Y(n974) );
  OAI2BB2XL U1898 ( .B0(n2039), .B1(n2141), .A0N(\register[28][29] ), .A1N(
        n2143), .Y(n975) );
  OAI2BB2XL U1899 ( .B0(n2036), .B1(n2141), .A0N(\register[28][30] ), .A1N(
        n2143), .Y(n976) );
  OAI2BB2XL U1900 ( .B0(n2033), .B1(n2141), .A0N(\register[28][31] ), .A1N(
        n2143), .Y(n977) );
  OAI2BB2XL U1901 ( .B0(n2126), .B1(n2137), .A0N(\register[29][0] ), .A1N(
        n2139), .Y(n978) );
  OAI2BB2XL U1902 ( .B0(n2123), .B1(n2137), .A0N(\register[29][1] ), .A1N(
        n2140), .Y(n979) );
  OAI2BB2XL U1903 ( .B0(n2120), .B1(n2137), .A0N(\register[29][2] ), .A1N(
        n2140), .Y(n980) );
  OAI2BB2XL U1904 ( .B0(n2117), .B1(n2137), .A0N(\register[29][3] ), .A1N(
        n2140), .Y(n981) );
  OAI2BB2XL U1905 ( .B0(n2114), .B1(n2137), .A0N(\register[29][4] ), .A1N(
        n2140), .Y(n982) );
  OAI2BB2XL U1906 ( .B0(n2111), .B1(n2137), .A0N(\register[29][5] ), .A1N(
        n2140), .Y(n983) );
  OAI2BB2XL U1907 ( .B0(n2108), .B1(n2137), .A0N(\register[29][6] ), .A1N(
        n2140), .Y(n984) );
  OAI2BB2XL U1908 ( .B0(n2105), .B1(n2137), .A0N(\register[29][7] ), .A1N(
        n2140), .Y(n985) );
  OAI2BB2XL U1909 ( .B0(n2102), .B1(n2138), .A0N(\register[29][8] ), .A1N(
        n2140), .Y(n986) );
  OAI2BB2XL U1910 ( .B0(n2099), .B1(n2138), .A0N(\register[29][9] ), .A1N(
        n2140), .Y(n987) );
  OAI2BB2XL U1911 ( .B0(n2096), .B1(n2138), .A0N(\register[29][10] ), .A1N(
        n2140), .Y(n988) );
  OAI2BB2XL U1912 ( .B0(n2093), .B1(n2138), .A0N(\register[29][11] ), .A1N(
        n2140), .Y(n989) );
  OAI2BB2XL U1913 ( .B0(n2090), .B1(n2138), .A0N(\register[29][12] ), .A1N(
        n2140), .Y(n990) );
  OAI2BB2XL U1914 ( .B0(n2087), .B1(n2138), .A0N(\register[29][13] ), .A1N(
        n2140), .Y(n991) );
  OAI2BB2XL U1915 ( .B0(n2084), .B1(n2138), .A0N(\register[29][14] ), .A1N(
        n2140), .Y(n992) );
  OAI2BB2XL U1916 ( .B0(n2081), .B1(n2138), .A0N(\register[29][15] ), .A1N(
        n2140), .Y(n993) );
  OAI2BB2XL U1917 ( .B0(n2078), .B1(n2139), .A0N(\register[29][16] ), .A1N(
        n2140), .Y(n994) );
  OAI2BB2XL U1918 ( .B0(n2075), .B1(n2139), .A0N(\register[29][17] ), .A1N(
        n2140), .Y(n995) );
  OAI2BB2XL U1919 ( .B0(n2072), .B1(n2138), .A0N(\register[29][18] ), .A1N(
        n2140), .Y(n996) );
  OAI2BB2XL U1920 ( .B0(n2069), .B1(n2139), .A0N(\register[29][19] ), .A1N(
        n2140), .Y(n997) );
  OAI2BB2XL U1921 ( .B0(n2066), .B1(n2139), .A0N(\register[29][20] ), .A1N(
        n2140), .Y(n998) );
  OAI2BB2XL U1922 ( .B0(n2063), .B1(n2139), .A0N(\register[29][21] ), .A1N(
        n2139), .Y(n999) );
  OAI2BB2XL U1923 ( .B0(n2060), .B1(n2139), .A0N(\register[29][22] ), .A1N(
        n2139), .Y(n1000) );
  OAI2BB2XL U1924 ( .B0(n2057), .B1(n2139), .A0N(\register[29][23] ), .A1N(
        n2139), .Y(n1001) );
  OAI2BB2XL U1925 ( .B0(n2054), .B1(n2139), .A0N(\register[29][24] ), .A1N(
        n2139), .Y(n1002) );
  OAI2BB2XL U1926 ( .B0(n2051), .B1(n2138), .A0N(\register[29][25] ), .A1N(
        n2139), .Y(n1003) );
  OAI2BB2XL U1927 ( .B0(n2048), .B1(n2138), .A0N(\register[29][26] ), .A1N(
        n2139), .Y(n1004) );
  OAI2BB2XL U1928 ( .B0(n2045), .B1(n2138), .A0N(\register[29][27] ), .A1N(
        n2139), .Y(n1005) );
  OAI2BB2XL U1929 ( .B0(n2042), .B1(n2137), .A0N(\register[29][28] ), .A1N(
        n2139), .Y(n1006) );
  OAI2BB2XL U1930 ( .B0(n2039), .B1(n2137), .A0N(\register[29][29] ), .A1N(
        n2139), .Y(n1007) );
  OAI2BB2XL U1931 ( .B0(n2036), .B1(n2137), .A0N(\register[29][30] ), .A1N(
        n2139), .Y(n1008) );
  OAI2BB2XL U1932 ( .B0(n2033), .B1(n2137), .A0N(\register[29][31] ), .A1N(
        n2139), .Y(n1009) );
  OAI2BB2XL U1933 ( .B0(n2126), .B1(n2133), .A0N(\register[30][0] ), .A1N(
        n2135), .Y(n1010) );
  OAI2BB2XL U1934 ( .B0(n2123), .B1(n2133), .A0N(\register[30][1] ), .A1N(
        n2136), .Y(n1011) );
  OAI2BB2XL U1935 ( .B0(n2120), .B1(n2133), .A0N(\register[30][2] ), .A1N(
        n2136), .Y(n1012) );
  OAI2BB2XL U1936 ( .B0(n2117), .B1(n2133), .A0N(\register[30][3] ), .A1N(
        n2136), .Y(n1013) );
  OAI2BB2XL U1937 ( .B0(n2114), .B1(n2133), .A0N(\register[30][4] ), .A1N(
        n2136), .Y(n1014) );
  OAI2BB2XL U1938 ( .B0(n2111), .B1(n2133), .A0N(\register[30][5] ), .A1N(
        n2136), .Y(n1015) );
  OAI2BB2XL U1939 ( .B0(n2108), .B1(n2133), .A0N(\register[30][6] ), .A1N(
        n2136), .Y(n1016) );
  OAI2BB2XL U1940 ( .B0(n2105), .B1(n2133), .A0N(\register[30][7] ), .A1N(
        n2136), .Y(n1017) );
  OAI2BB2XL U1941 ( .B0(n2102), .B1(n2134), .A0N(\register[30][8] ), .A1N(
        n2136), .Y(n1018) );
  OAI2BB2XL U1942 ( .B0(n2099), .B1(n2134), .A0N(\register[30][9] ), .A1N(
        n2136), .Y(n1019) );
  OAI2BB2XL U1943 ( .B0(n2096), .B1(n2134), .A0N(\register[30][10] ), .A1N(
        n2136), .Y(n1020) );
  OAI2BB2XL U1944 ( .B0(n2093), .B1(n2134), .A0N(\register[30][11] ), .A1N(
        n2136), .Y(n1021) );
  OAI2BB2XL U1945 ( .B0(n2090), .B1(n2134), .A0N(\register[30][12] ), .A1N(
        n2136), .Y(n1022) );
  OAI2BB2XL U1946 ( .B0(n2087), .B1(n2134), .A0N(\register[30][13] ), .A1N(
        n2136), .Y(n1023) );
  OAI2BB2XL U1947 ( .B0(n2084), .B1(n2134), .A0N(\register[30][14] ), .A1N(
        n2136), .Y(n1024) );
  OAI2BB2XL U1948 ( .B0(n2081), .B1(n2134), .A0N(\register[30][15] ), .A1N(
        n2136), .Y(n1025) );
  OAI2BB2XL U1949 ( .B0(n2078), .B1(n2135), .A0N(\register[30][16] ), .A1N(
        n2136), .Y(n1026) );
  OAI2BB2XL U1950 ( .B0(n2075), .B1(n2135), .A0N(\register[30][17] ), .A1N(
        n2136), .Y(n1027) );
  OAI2BB2XL U1951 ( .B0(n2072), .B1(n2134), .A0N(\register[30][18] ), .A1N(
        n2136), .Y(n1028) );
  OAI2BB2XL U1952 ( .B0(n2069), .B1(n2135), .A0N(\register[30][19] ), .A1N(
        n2136), .Y(n1029) );
  OAI2BB2XL U1953 ( .B0(n2066), .B1(n2135), .A0N(\register[30][20] ), .A1N(
        n2136), .Y(n1030) );
  OAI2BB2XL U1954 ( .B0(n2063), .B1(n2135), .A0N(\register[30][21] ), .A1N(
        n2135), .Y(n1031) );
  OAI2BB2XL U1955 ( .B0(n2060), .B1(n2135), .A0N(\register[30][22] ), .A1N(
        n2135), .Y(n1032) );
  OAI2BB2XL U1956 ( .B0(n2057), .B1(n2135), .A0N(\register[30][23] ), .A1N(
        n2135), .Y(n1033) );
  OAI2BB2XL U1957 ( .B0(n2054), .B1(n2135), .A0N(\register[30][24] ), .A1N(
        n2135), .Y(n1034) );
  OAI2BB2XL U1958 ( .B0(n2051), .B1(n2134), .A0N(\register[30][25] ), .A1N(
        n2135), .Y(n1035) );
  OAI2BB2XL U1959 ( .B0(n2048), .B1(n2134), .A0N(\register[30][26] ), .A1N(
        n2135), .Y(n1036) );
  OAI2BB2XL U1960 ( .B0(n2045), .B1(n2134), .A0N(\register[30][27] ), .A1N(
        n2135), .Y(n1037) );
  OAI2BB2XL U1961 ( .B0(n2042), .B1(n2133), .A0N(\register[30][28] ), .A1N(
        n2135), .Y(n1038) );
  OAI2BB2XL U1962 ( .B0(n2039), .B1(n2133), .A0N(\register[30][29] ), .A1N(
        n2135), .Y(n1039) );
  OAI2BB2XL U1963 ( .B0(n2036), .B1(n2133), .A0N(\register[30][30] ), .A1N(
        n2135), .Y(n1040) );
  OAI2BB2XL U1964 ( .B0(n2033), .B1(n2133), .A0N(\register[30][31] ), .A1N(
        n2135), .Y(n1041) );
  OAI2BB2XL U1965 ( .B0(n2126), .B1(n2129), .A0N(\register[31][0] ), .A1N(
        n2131), .Y(n1042) );
  OAI2BB2XL U1966 ( .B0(n2123), .B1(n2129), .A0N(\register[31][1] ), .A1N(
        n2132), .Y(n1043) );
  OAI2BB2XL U1967 ( .B0(n2120), .B1(n2129), .A0N(\register[31][2] ), .A1N(
        n2132), .Y(n1044) );
  OAI2BB2XL U1968 ( .B0(n2117), .B1(n2129), .A0N(\register[31][3] ), .A1N(
        n2132), .Y(n1045) );
  OAI2BB2XL U1969 ( .B0(n2114), .B1(n2129), .A0N(\register[31][4] ), .A1N(
        n2132), .Y(n1046) );
  OAI2BB2XL U1970 ( .B0(n2111), .B1(n2129), .A0N(\register[31][5] ), .A1N(
        n2132), .Y(n1047) );
  OAI2BB2XL U1971 ( .B0(n2108), .B1(n2129), .A0N(\register[31][6] ), .A1N(
        n2132), .Y(n1048) );
  OAI2BB2XL U1972 ( .B0(n2105), .B1(n2129), .A0N(\register[31][7] ), .A1N(
        n2132), .Y(n1049) );
  OAI2BB2XL U1973 ( .B0(n2102), .B1(n2130), .A0N(\register[31][8] ), .A1N(
        n2132), .Y(n1050) );
  OAI2BB2XL U1974 ( .B0(n2099), .B1(n2130), .A0N(\register[31][9] ), .A1N(
        n2132), .Y(n1051) );
  OAI2BB2XL U1975 ( .B0(n2096), .B1(n2130), .A0N(\register[31][10] ), .A1N(
        n2132), .Y(n1052) );
  OAI2BB2XL U1976 ( .B0(n2093), .B1(n2130), .A0N(\register[31][11] ), .A1N(
        n2132), .Y(n1053) );
  OAI2BB2XL U1977 ( .B0(n2090), .B1(n2130), .A0N(\register[31][12] ), .A1N(
        n2132), .Y(n1054) );
  OAI2BB2XL U1978 ( .B0(n2087), .B1(n2130), .A0N(\register[31][13] ), .A1N(
        n2132), .Y(n1055) );
  OAI2BB2XL U1979 ( .B0(n2084), .B1(n2130), .A0N(\register[31][14] ), .A1N(
        n2132), .Y(n1056) );
  OAI2BB2XL U1980 ( .B0(n2081), .B1(n2130), .A0N(\register[31][15] ), .A1N(
        n2132), .Y(n1057) );
  OAI2BB2XL U1981 ( .B0(n2078), .B1(n2131), .A0N(\register[31][16] ), .A1N(
        n2132), .Y(n1058) );
  OAI2BB2XL U1982 ( .B0(n2075), .B1(n2131), .A0N(\register[31][17] ), .A1N(
        n2132), .Y(n1059) );
  OAI2BB2XL U1983 ( .B0(n2072), .B1(n2130), .A0N(\register[31][18] ), .A1N(
        n2132), .Y(n1060) );
  OAI2BB2XL U1984 ( .B0(n2069), .B1(n2131), .A0N(\register[31][19] ), .A1N(
        n2132), .Y(n1061) );
  OAI2BB2XL U1985 ( .B0(n2066), .B1(n2131), .A0N(\register[31][20] ), .A1N(
        n2132), .Y(n1062) );
  OAI2BB2XL U1986 ( .B0(n2063), .B1(n2131), .A0N(\register[31][21] ), .A1N(
        n2131), .Y(n1063) );
  OAI2BB2XL U1987 ( .B0(n2060), .B1(n2131), .A0N(\register[31][22] ), .A1N(
        n2131), .Y(n1064) );
  OAI2BB2XL U1988 ( .B0(n2057), .B1(n2131), .A0N(\register[31][23] ), .A1N(
        n2131), .Y(n1065) );
  OAI2BB2XL U1989 ( .B0(n2054), .B1(n2131), .A0N(\register[31][24] ), .A1N(
        n2131), .Y(n1066) );
  OAI2BB2XL U1990 ( .B0(n2051), .B1(n2130), .A0N(\register[31][25] ), .A1N(
        n2131), .Y(n1067) );
  OAI2BB2XL U1991 ( .B0(n2048), .B1(n2130), .A0N(\register[31][26] ), .A1N(
        n2131), .Y(n1068) );
  OAI2BB2XL U1992 ( .B0(n2045), .B1(n2130), .A0N(\register[31][27] ), .A1N(
        n2131), .Y(n1069) );
  OAI2BB2XL U1993 ( .B0(n2042), .B1(n2129), .A0N(\register[31][28] ), .A1N(
        n2131), .Y(n1070) );
  OAI2BB2XL U1994 ( .B0(n2039), .B1(n2129), .A0N(\register[31][29] ), .A1N(
        n2131), .Y(n1071) );
  OAI2BB2XL U1995 ( .B0(n2036), .B1(n2129), .A0N(\register[31][30] ), .A1N(
        n2131), .Y(n1072) );
  OAI2BB2XL U1996 ( .B0(n2033), .B1(n2129), .A0N(\register[31][31] ), .A1N(
        n2131), .Y(n1073) );
  OAI2BB2XL U1997 ( .B0(n2249), .B1(n2128), .A0N(\register[1][0] ), .A1N(n2251), .Y(n82) );
  OAI2BB2XL U1998 ( .B0(n2249), .B1(n2125), .A0N(\register[1][1] ), .A1N(n2252), .Y(n83) );
  OAI2BB2XL U1999 ( .B0(n2249), .B1(n2122), .A0N(\register[1][2] ), .A1N(n2252), .Y(n84) );
  OAI2BB2XL U2000 ( .B0(n2249), .B1(n2119), .A0N(\register[1][3] ), .A1N(n2252), .Y(n85) );
  OAI2BB2XL U2001 ( .B0(n2249), .B1(n2116), .A0N(\register[1][4] ), .A1N(n2252), .Y(n86) );
  OAI2BB2XL U2002 ( .B0(n2249), .B1(n2113), .A0N(\register[1][5] ), .A1N(n2252), .Y(n87) );
  OAI2BB2XL U2003 ( .B0(n2249), .B1(n2110), .A0N(\register[1][6] ), .A1N(n2252), .Y(n88) );
  OAI2BB2XL U2004 ( .B0(n2249), .B1(n2107), .A0N(\register[1][7] ), .A1N(n2252), .Y(n89) );
  OAI2BB2XL U2005 ( .B0(n2250), .B1(n2104), .A0N(\register[1][8] ), .A1N(n2252), .Y(n90) );
  OAI2BB2XL U2006 ( .B0(n2250), .B1(n2101), .A0N(\register[1][9] ), .A1N(n2252), .Y(n91) );
  OAI2BB2XL U2007 ( .B0(n2250), .B1(n2098), .A0N(\register[1][10] ), .A1N(
        n2252), .Y(n92) );
  OAI2BB2XL U2008 ( .B0(n2250), .B1(n2095), .A0N(\register[1][11] ), .A1N(
        n2252), .Y(n93) );
  OAI2BB2XL U2009 ( .B0(n2250), .B1(n2092), .A0N(\register[1][12] ), .A1N(
        n2252), .Y(n94) );
  OAI2BB2XL U2010 ( .B0(n2250), .B1(n2089), .A0N(\register[1][13] ), .A1N(
        n2252), .Y(n95) );
  OAI2BB2XL U2011 ( .B0(n2250), .B1(n2086), .A0N(\register[1][14] ), .A1N(
        n2252), .Y(n96) );
  OAI2BB2XL U2012 ( .B0(n2250), .B1(n2083), .A0N(\register[1][15] ), .A1N(
        n2252), .Y(n97) );
  OAI2BB2XL U2013 ( .B0(n2251), .B1(n2080), .A0N(\register[1][16] ), .A1N(
        n2252), .Y(n98) );
  OAI2BB2XL U2014 ( .B0(n2251), .B1(n2077), .A0N(\register[1][17] ), .A1N(
        n2252), .Y(n99) );
  OAI2BB2XL U2015 ( .B0(n2250), .B1(n2074), .A0N(\register[1][18] ), .A1N(
        n2252), .Y(n100) );
  OAI2BB2XL U2016 ( .B0(n2251), .B1(n2071), .A0N(\register[1][19] ), .A1N(
        n2252), .Y(n101) );
  OAI2BB2XL U2017 ( .B0(n2251), .B1(n2068), .A0N(\register[1][20] ), .A1N(
        n2251), .Y(n102) );
  OAI2BB2XL U2018 ( .B0(n2251), .B1(n2065), .A0N(\register[1][21] ), .A1N(
        n2251), .Y(n103) );
  OAI2BB2XL U2019 ( .B0(n2251), .B1(n2062), .A0N(\register[1][22] ), .A1N(
        n2251), .Y(n104) );
  OAI2BB2XL U2020 ( .B0(n2251), .B1(n2059), .A0N(\register[1][23] ), .A1N(
        n2251), .Y(n105) );
  OAI2BB2XL U2021 ( .B0(n2251), .B1(n2056), .A0N(\register[1][24] ), .A1N(
        n2251), .Y(n106) );
  OAI2BB2XL U2022 ( .B0(n2250), .B1(n2053), .A0N(\register[1][25] ), .A1N(
        n2251), .Y(n107) );
  OAI2BB2XL U2023 ( .B0(n2250), .B1(n2050), .A0N(\register[1][26] ), .A1N(
        n2251), .Y(n108) );
  OAI2BB2XL U2024 ( .B0(n2250), .B1(n2047), .A0N(\register[1][27] ), .A1N(
        n2251), .Y(n109) );
  OAI2BB2XL U2025 ( .B0(n2249), .B1(n2044), .A0N(\register[1][28] ), .A1N(
        n2251), .Y(n110) );
  OAI2BB2XL U2026 ( .B0(n2249), .B1(n2041), .A0N(\register[1][29] ), .A1N(
        n2251), .Y(n111) );
  OAI2BB2XL U2027 ( .B0(n2249), .B1(n2038), .A0N(\register[1][30] ), .A1N(
        n2251), .Y(n112) );
  OAI2BB2XL U2028 ( .B0(n2249), .B1(n2035), .A0N(\register[1][31] ), .A1N(
        n2251), .Y(n113) );
  NAND2BX1 U2029 ( .AN(n1424), .B(n1423), .Y(n1190) );
  OAI22XL U2030 ( .A0(n1495), .A1(n1524), .B0(n1492), .B1(\register[1][10] ), 
        .Y(n1424) );
  NAND2BX1 U2031 ( .AN(n1427), .B(n1426), .Y(n1182) );
  OAI22XL U2032 ( .A0(n1495), .A1(n1524), .B0(n1492), .B1(\register[1][9] ), 
        .Y(n1427) );
  NAND2BX1 U2033 ( .AN(n1421), .B(n1420), .Y(n1198) );
  OAI22XL U2034 ( .A0(n1494), .A1(n1524), .B0(n1492), .B1(\register[1][11] ), 
        .Y(n1421) );
  NAND2BX1 U2035 ( .AN(n1418), .B(n1417), .Y(n1206) );
  OAI22XL U2036 ( .A0(n1494), .A1(n1524), .B0(n1493), .B1(\register[1][12] ), 
        .Y(n1418) );
  NAND2BX1 U2037 ( .AN(n1415), .B(n1414), .Y(n1214) );
  OAI22XL U2038 ( .A0(n1494), .A1(n1525), .B0(n1492), .B1(\register[1][13] ), 
        .Y(n1415) );
  NAND2BX1 U2039 ( .AN(n1412), .B(n1411), .Y(n1222) );
  MXI2X1 U2040 ( .A(n2379), .B(n1410), .S0(n1527), .Y(n1411) );
  OAI22XL U2041 ( .A0(n1495), .A1(n1525), .B0(n1492), .B1(\register[1][14] ), 
        .Y(n1412) );
  NAND2BX1 U2042 ( .AN(n1403), .B(n1402), .Y(n1246) );
  MXI2X1 U2043 ( .A(n2382), .B(n1401), .S0(n1527), .Y(n1402) );
  OAI22XL U2044 ( .A0(n1494), .A1(n1525), .B0(n1493), .B1(\register[1][17] ), 
        .Y(n1403) );
  NOR2BX1 U2045 ( .AN(n1491), .B(\register[3][17] ), .Y(n1401) );
  NAND2BX1 U2046 ( .AN(n1909), .B(n1908), .Y(n1719) );
  MXI2X1 U2047 ( .A(n2379), .B(n1907), .S0(n2024), .Y(n1908) );
  OAI22XL U2048 ( .A0(n1992), .A1(n2022), .B0(n1989), .B1(\register[1][14] ), 
        .Y(n1909) );
  NOR2BX1 U2049 ( .AN(n1988), .B(\register[3][14] ), .Y(n1907) );
  NAND2BX1 U2050 ( .AN(n1900), .B(n1899), .Y(n1743) );
  MXI2X1 U2051 ( .A(n2382), .B(n1898), .S0(n2024), .Y(n1899) );
  OAI22XL U2052 ( .A0(n1991), .A1(n2022), .B0(n1990), .B1(\register[1][17] ), 
        .Y(n1900) );
  NOR2BX1 U2053 ( .AN(n1988), .B(\register[3][17] ), .Y(n1898) );
  NAND2BX1 U2054 ( .AN(n1882), .B(n1881), .Y(n1791) );
  MXI2X1 U2055 ( .A(n2388), .B(n1880), .S0(n2024), .Y(n1881) );
  OAI22XL U2056 ( .A0(n1992), .A1(n2022), .B0(n1990), .B1(\register[1][23] ), 
        .Y(n1882) );
  NOR2BX1 U2057 ( .AN(n1988), .B(\register[3][23] ), .Y(n1880) );
  NAND2BX1 U2058 ( .AN(n1876), .B(n1875), .Y(n1807) );
  MXI2X1 U2059 ( .A(n2390), .B(n1874), .S0(n2024), .Y(n1875) );
  OAI22XL U2060 ( .A0(n1992), .A1(n2022), .B0(n1991), .B1(\register[1][25] ), 
        .Y(n1876) );
  NOR2BX1 U2061 ( .AN(n1988), .B(\register[3][25] ), .Y(n1874) );
  NAND2BX1 U2062 ( .AN(n1873), .B(n1872), .Y(n1815) );
  MXI2X1 U2063 ( .A(n2391), .B(n1871), .S0(n2024), .Y(n1872) );
  OAI22XL U2064 ( .A0(n1992), .A1(n2023), .B0(n1990), .B1(\register[1][26] ), 
        .Y(n1873) );
  NOR2BX1 U2065 ( .AN(n1988), .B(\register[3][26] ), .Y(n1871) );
  NAND2BX1 U2066 ( .AN(n1870), .B(n1869), .Y(n1823) );
  MXI2X1 U2067 ( .A(n2392), .B(n1868), .S0(n2024), .Y(n1869) );
  OAI22XL U2068 ( .A0(n1993), .A1(n2023), .B0(n1991), .B1(\register[1][27] ), 
        .Y(n1870) );
  NOR2BX1 U2069 ( .AN(n1988), .B(\register[3][27] ), .Y(n1868) );
  NAND2BX1 U2070 ( .AN(n1867), .B(n1866), .Y(n1831) );
  MXI2X1 U2071 ( .A(n2393), .B(n1865), .S0(n2025), .Y(n1866) );
  OAI22XL U2072 ( .A0(n1993), .A1(n2022), .B0(n1991), .B1(\register[1][28] ), 
        .Y(n1867) );
  NOR2BX1 U2073 ( .AN(n1988), .B(\register[3][28] ), .Y(n1865) );
  NAND2BX1 U2074 ( .AN(n1864), .B(n1863), .Y(n1839) );
  MXI2X1 U2075 ( .A(n2394), .B(n1862), .S0(n2025), .Y(n1863) );
  OAI22XL U2076 ( .A0(n1993), .A1(n2023), .B0(n1991), .B1(\register[1][29] ), 
        .Y(n1864) );
  NOR2BX1 U2077 ( .AN(n1988), .B(\register[3][29] ), .Y(n1862) );
  NAND2BX1 U2078 ( .AN(n1861), .B(n1860), .Y(n1847) );
  MXI2X1 U2079 ( .A(n2395), .B(n1859), .S0(n2025), .Y(n1860) );
  OAI22XL U2080 ( .A0(n1993), .A1(n2023), .B0(n1990), .B1(\register[1][30] ), 
        .Y(n1861) );
  NOR2BX1 U2081 ( .AN(n1988), .B(\register[3][30] ), .Y(n1859) );
  NAND2BX1 U2082 ( .AN(n1858), .B(n1857), .Y(n1855) );
  MXI2X1 U2083 ( .A(n2396), .B(n1856), .S0(n2025), .Y(n1857) );
  OAI22XL U2084 ( .A0(n1993), .A1(n2022), .B0(n1991), .B1(\register[1][31] ), 
        .Y(n1858) );
  NOR2BX1 U2085 ( .AN(n1988), .B(\register[3][31] ), .Y(n1856) );
  NAND2BX1 U2086 ( .AN(n1409), .B(n1408), .Y(n1230) );
  MXI2X1 U2087 ( .A(n2380), .B(n1407), .S0(n1526), .Y(n1408) );
  OAI22XL U2088 ( .A0(n1494), .A1(n1525), .B0(n1493), .B1(\register[1][15] ), 
        .Y(n1409) );
  NOR2BX1 U2089 ( .AN(n1491), .B(\register[3][15] ), .Y(n1407) );
  NAND2BX1 U2090 ( .AN(n1406), .B(n1405), .Y(n1238) );
  MXI2X1 U2091 ( .A(n2381), .B(n1404), .S0(n1526), .Y(n1405) );
  OAI22XL U2092 ( .A0(n1495), .A1(n1525), .B0(n1493), .B1(\register[1][16] ), 
        .Y(n1406) );
  NOR2BX1 U2093 ( .AN(n1491), .B(\register[3][16] ), .Y(n1404) );
  NAND2BX1 U2094 ( .AN(n1400), .B(n1399), .Y(n1254) );
  MXI2X1 U2095 ( .A(n2383), .B(n1398), .S0(n1526), .Y(n1399) );
  OAI22XL U2096 ( .A0(n1494), .A1(n1525), .B0(n1493), .B1(\register[1][18] ), 
        .Y(n1400) );
  NOR2BX1 U2097 ( .AN(n1491), .B(\register[3][18] ), .Y(n1398) );
  NAND2BX1 U2098 ( .AN(n1397), .B(n1396), .Y(n1262) );
  MXI2X1 U2099 ( .A(n2384), .B(n1395), .S0(n1526), .Y(n1396) );
  OAI22XL U2100 ( .A0(n1494), .A1(n1525), .B0(n1493), .B1(\register[1][19] ), 
        .Y(n1397) );
  NOR2BX1 U2101 ( .AN(n1491), .B(\register[3][19] ), .Y(n1395) );
  NAND2BX1 U2102 ( .AN(n1394), .B(n1393), .Y(n1270) );
  MXI2X1 U2103 ( .A(n2385), .B(n1392), .S0(n1526), .Y(n1393) );
  OAI22XL U2104 ( .A0(n1495), .A1(n1525), .B0(n1493), .B1(\register[1][20] ), 
        .Y(n1394) );
  NOR2BX1 U2105 ( .AN(n1491), .B(\register[3][20] ), .Y(n1392) );
  NAND2BX1 U2106 ( .AN(n1391), .B(n1390), .Y(n1278) );
  MXI2X1 U2107 ( .A(n2386), .B(n1389), .S0(n1526), .Y(n1390) );
  OAI22XL U2108 ( .A0(n1494), .A1(n1525), .B0(n1493), .B1(\register[1][21] ), 
        .Y(n1391) );
  NOR2BX1 U2109 ( .AN(n1491), .B(\register[3][21] ), .Y(n1389) );
  NAND2BX1 U2110 ( .AN(n1388), .B(n1387), .Y(n1286) );
  MXI2X1 U2111 ( .A(n2387), .B(n1386), .S0(n1526), .Y(n1387) );
  OAI22XL U2112 ( .A0(n1495), .A1(n1525), .B0(n1493), .B1(\register[1][22] ), 
        .Y(n1388) );
  NOR2BX1 U2113 ( .AN(n1491), .B(\register[3][22] ), .Y(n1386) );
  NAND2BX1 U2114 ( .AN(n1906), .B(n1905), .Y(n1727) );
  MXI2X1 U2115 ( .A(n2380), .B(n1904), .S0(n2023), .Y(n1905) );
  OAI22XL U2116 ( .A0(n1991), .A1(n2022), .B0(n1990), .B1(\register[1][15] ), 
        .Y(n1906) );
  NOR2BX1 U2117 ( .AN(n1988), .B(\register[3][15] ), .Y(n1904) );
  NAND2BX1 U2118 ( .AN(n1903), .B(n1902), .Y(n1735) );
  MXI2X1 U2119 ( .A(n2381), .B(n1901), .S0(n2023), .Y(n1902) );
  OAI22XL U2120 ( .A0(n1992), .A1(n2022), .B0(n1990), .B1(\register[1][16] ), 
        .Y(n1903) );
  NOR2BX1 U2121 ( .AN(n1988), .B(\register[3][16] ), .Y(n1901) );
  NAND2BX1 U2122 ( .AN(n1897), .B(n1896), .Y(n1751) );
  MXI2X1 U2123 ( .A(n2383), .B(n1895), .S0(n2023), .Y(n1896) );
  OAI22XL U2124 ( .A0(n1991), .A1(n2022), .B0(n1990), .B1(\register[1][18] ), 
        .Y(n1897) );
  NOR2BX1 U2125 ( .AN(n1988), .B(\register[3][18] ), .Y(n1895) );
  NAND2BX1 U2126 ( .AN(n1894), .B(n1893), .Y(n1759) );
  MXI2X1 U2127 ( .A(n2384), .B(n1892), .S0(n2023), .Y(n1893) );
  OAI22XL U2128 ( .A0(n1991), .A1(n2022), .B0(n1990), .B1(\register[1][19] ), 
        .Y(n1894) );
  NOR2BX1 U2129 ( .AN(n1988), .B(\register[3][19] ), .Y(n1892) );
  NAND2BX1 U2130 ( .AN(n1891), .B(n1890), .Y(n1767) );
  MXI2X1 U2131 ( .A(n2385), .B(n1889), .S0(n2023), .Y(n1890) );
  OAI22XL U2132 ( .A0(n1992), .A1(n2022), .B0(n1990), .B1(\register[1][20] ), 
        .Y(n1891) );
  NOR2BX1 U2133 ( .AN(n1988), .B(\register[3][20] ), .Y(n1889) );
  NAND2BX1 U2134 ( .AN(n1888), .B(n1887), .Y(n1775) );
  MXI2X1 U2135 ( .A(n2386), .B(n1886), .S0(n2023), .Y(n1887) );
  OAI22XL U2136 ( .A0(n1991), .A1(n2022), .B0(n1990), .B1(\register[1][21] ), 
        .Y(n1888) );
  NOR2BX1 U2137 ( .AN(n1988), .B(\register[3][21] ), .Y(n1886) );
  NAND2BX1 U2138 ( .AN(n1885), .B(n1884), .Y(n1783) );
  MXI2X1 U2139 ( .A(n2387), .B(n1883), .S0(n2023), .Y(n1884) );
  OAI22XL U2140 ( .A0(n1992), .A1(n2022), .B0(n1990), .B1(\register[1][22] ), 
        .Y(n1885) );
  NOR2BX1 U2141 ( .AN(n1988), .B(\register[3][22] ), .Y(n1883) );
  NAND2BX1 U2142 ( .AN(n1879), .B(n1878), .Y(n1799) );
  MXI2X1 U2143 ( .A(n2389), .B(n1877), .S0(n2023), .Y(n1878) );
  OAI22XL U2144 ( .A0(n1993), .A1(n2023), .B0(n1990), .B1(\register[1][24] ), 
        .Y(n1879) );
  NOR2BX1 U2145 ( .AN(n1988), .B(\register[3][24] ), .Y(n1877) );
  MXI4X1 U2146 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1520), .S1(n1489), .Y(
        n1229) );
  MXI4X1 U2147 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1523), .S1(n1489), 
        .Y(n1225) );
  MXI4X1 U2148 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1511), .S1(n1485), .Y(
        n1245) );
  MXI4X1 U2149 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1241) );
  MXI4X1 U2150 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1512), .S1(n1485), .Y(
        n1253) );
  MXI4X1 U2151 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1511), .S1(n1485), 
        .Y(n1249) );
  MXI4X1 U2152 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1512), .S1(n1485), .Y(
        n1261) );
  MXI4X1 U2153 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1257) );
  MXI4X1 U2154 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1513), .S1(n1485), .Y(
        n1269) );
  MXI4X1 U2155 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1265) );
  MXI4X1 U2156 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1513), .S1(n1486), .Y(
        n1277) );
  MXI4X1 U2157 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1513), .S1(n1485), 
        .Y(n1273) );
  MXI4X1 U2158 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1513), .S1(n1486), .Y(
        n1285) );
  MXI4X1 U2159 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1281) );
  MXI4X1 U2160 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n2018), .S1(n1987), .Y(
        n1674) );
  MXI4X1 U2161 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n2018), .S1(n1987), .Y(
        n1678) );
  MXI4X1 U2162 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n2018), .S1(n1987), 
        .Y(n1682) );
  MXI4X1 U2163 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n2019), .S1(n1987), .Y(
        n1686) );
  MXI4X1 U2164 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1690) );
  MXI4X1 U2165 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n2019), .S1(n1987), .Y(
        n1694) );
  MXI4X1 U2166 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1698) );
  MXI4X1 U2167 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n2019), .S1(n1987), .Y(
        n1702) );
  MXI4X1 U2168 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n2020), .S1(n1986), 
        .Y(n1706) );
  MXI4X1 U2169 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n2020), .S1(n1986), .Y(
        n1710) );
  MXI4X1 U2170 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n2020), .S1(n1986), .Y(
        n1718) );
  MXI4X1 U2171 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1714) );
  MXI4X1 U2172 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n2017), .S1(n1986), .Y(
        n1726) );
  MXI4X1 U2173 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n2020), .S1(n1986), 
        .Y(n1722) );
  MXI4X1 U2174 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n2008), .S1(n1982), .Y(
        n1734) );
  MXI4X1 U2175 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n2008), .S1(n1981), 
        .Y(n1730) );
  MXI4X1 U2176 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n2008), .S1(n1982), .Y(
        n1742) );
  MXI4X1 U2177 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1738) );
  MXI4X1 U2178 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n2009), .S1(n1982), .Y(
        n1750) );
  MXI4X1 U2179 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n2008), .S1(n1982), 
        .Y(n1746) );
  MXI4X1 U2180 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n2009), .S1(n1982), .Y(
        n1758) );
  MXI4X1 U2181 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1754) );
  MXI4X1 U2182 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n2010), .S1(n1982), .Y(
        n1766) );
  MXI4X1 U2183 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1762) );
  MXI4X1 U2184 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n2010), .S1(n1983), .Y(
        n1774) );
  MXI4X1 U2185 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n2010), .S1(n1982), 
        .Y(n1770) );
  MXI4X1 U2186 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n2010), .S1(n1983), .Y(
        n1782) );
  MXI4X1 U2187 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1778) );
  MXI4X1 U2188 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n2011), .S1(n1983), .Y(
        n1790) );
  MXI4X1 U2189 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n2011), .S1(n1983), 
        .Y(n1786) );
  MXI4X1 U2190 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n2011), .S1(n1983), .Y(
        n1798) );
  MXI4X1 U2191 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1794) );
  MXI4X1 U2192 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n2012), .S1(n1983), .Y(
        n1806) );
  MXI4X1 U2193 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n2011), .S1(n1983), 
        .Y(n1802) );
  MXI4X1 U2194 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n2012), .S1(n1984), .Y(
        n1814) );
  MXI4X1 U2195 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1810) );
  MXI4X1 U2196 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n2012), .S1(n1984), .Y(
        n1822) );
  MXI4X1 U2197 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1818) );
  MXI4X1 U2198 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n2013), .S1(n1984), .Y(
        n1830) );
  MXI4X1 U2199 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1826) );
  MXI4X1 U2200 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n2013), .S1(n1984), .Y(
        n1838) );
  MXI4X1 U2201 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1834) );
  MXI4X1 U2202 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n2014), .S1(n1984), .Y(
        n1846) );
  MXI4X1 U2203 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n2013), .S1(n1984), 
        .Y(n1842) );
  MXI4X1 U2204 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n2021), .S1(n1986), .Y(
        n1854) );
  MXI4X1 U2205 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n2014), .S1(n1984), 
        .Y(n1850) );
  MXI4X1 U2206 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1523), .S1(n1489), 
        .Y(n1226) );
  MXI4X1 U2207 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1242) );
  MXI4X1 U2208 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1512), .S1(n1485), 
        .Y(n1250) );
  MXI4X1 U2209 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1258) );
  MXI4X1 U2210 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1266) );
  MXI4X1 U2211 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1513), .S1(n1485), 
        .Y(n1274) );
  MXI4X1 U2212 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1282) );
  MXI4X1 U2213 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n2018), .S1(n1987), .Y(
        n1675) );
  MXI4X1 U2214 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n2018), .S1(n1987), 
        .Y(n1683) );
  MXI4X1 U2215 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1691) );
  MXI4X1 U2216 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1699) );
  MXI4X1 U2217 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n2020), .S1(n1986), 
        .Y(n1707) );
  MXI4X1 U2218 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1715) );
  MXI4X1 U2219 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n2020), .S1(n1986), 
        .Y(n1723) );
  MXI4X1 U2220 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n2008), .S1(n1982), 
        .Y(n1731) );
  MXI4X1 U2221 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1739) );
  MXI4X1 U2222 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n2009), .S1(n1982), 
        .Y(n1747) );
  MXI4X1 U2223 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1755) );
  MXI4X1 U2224 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1763) );
  MXI4X1 U2225 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n2010), .S1(n1982), 
        .Y(n1771) );
  MXI4X1 U2226 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1779) );
  MXI4X1 U2227 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n2011), .S1(n1983), 
        .Y(n1787) );
  MXI4X1 U2228 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1795) );
  MXI4X1 U2229 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n2011), .S1(n1983), 
        .Y(n1803) );
  MXI4X1 U2230 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1811) );
  MXI4X1 U2231 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1819) );
  MXI4X1 U2232 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1827) );
  MXI4X1 U2233 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1835) );
  MXI4X1 U2234 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n2014), .S1(n1984), 
        .Y(n1843) );
  MXI4X1 U2235 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n2014), .S1(n1984), 
        .Y(n1851) );
  MXI4X1 U2236 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1524), .S1(n1489), 
        .Y(n1227) );
  MXI4X1 U2237 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1243) );
  MXI4X1 U2238 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1512), .S1(n1485), 
        .Y(n1251) );
  MXI4X1 U2239 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1259) );
  MXI4X1 U2240 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1267) );
  MXI4X1 U2241 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1513), .S1(n1485), 
        .Y(n1275) );
  MXI4X1 U2242 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1283) );
  MXI4X1 U2243 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n2018), .S1(n1987), .Y(
        n1672) );
  MXI4X1 U2244 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n2018), .S1(n1987), .Y(
        n1676) );
  MXI4X1 U2245 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n2018), .S1(n1987), 
        .Y(n1680) );
  MXI4X1 U2246 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n2018), .S1(n1987), 
        .Y(n1684) );
  MXI4X1 U2247 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1688) );
  MXI4X1 U2248 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1692) );
  MXI4X1 U2249 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1696) );
  MXI4X1 U2250 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1700) );
  MXI4X1 U2251 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n2019), .S1(n1987), 
        .Y(n1704) );
  MXI4X1 U2252 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n2020), .S1(n1986), 
        .Y(n1708) );
  MXI4X1 U2253 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1716) );
  MXI4X1 U2254 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n2021), .S1(n1986), 
        .Y(n1724) );
  MXI4X1 U2255 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n2008), .S1(n1982), 
        .Y(n1732) );
  MXI4X1 U2256 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1740) );
  MXI4X1 U2257 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n2009), .S1(n1982), 
        .Y(n1748) );
  MXI4X1 U2258 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1756) );
  MXI4X1 U2259 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1764) );
  MXI4X1 U2260 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n2010), .S1(n1982), 
        .Y(n1772) );
  MXI4X1 U2261 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1780) );
  MXI4X1 U2262 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n2011), .S1(n1983), 
        .Y(n1788) );
  MXI4X1 U2263 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1796) );
  MXI4X1 U2264 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n2012), .S1(n1983), 
        .Y(n1804) );
  MXI4X1 U2265 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1812) );
  MXI4X1 U2266 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1820) );
  MXI4X1 U2267 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1828) );
  MXI4X1 U2268 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1836) );
  MXI4X1 U2269 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n2014), .S1(n1984), 
        .Y(n1844) );
  MXI4X1 U2270 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n2014), .S1(n1984), 
        .Y(n1852) );
  MXI4X1 U2271 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1524), .S1(n1489), 
        .Y(n1228) );
  MXI4X1 U2272 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1523), .S1(n1489), 
        .Y(n1224) );
  MXI4X1 U2273 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1244) );
  MXI4X1 U2274 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1511), .S1(n1485), 
        .Y(n1240) );
  MXI4X1 U2275 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1512), .S1(n1485), 
        .Y(n1252) );
  MXI4X1 U2276 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1511), .S1(n1485), 
        .Y(n1248) );
  MXI4X1 U2277 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1260) );
  MXI4X1 U2278 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1512), .S1(n1485), 
        .Y(n1256) );
  MXI4X1 U2279 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1268) );
  MXI4X1 U2280 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1512), .S1(n1485), 
        .Y(n1264) );
  MXI4X1 U2281 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1513), .S1(n1486), 
        .Y(n1276) );
  MXI4X1 U2282 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1513), .S1(n1485), 
        .Y(n1272) );
  MXI4X1 U2283 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1284) );
  MXI4X1 U2284 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1513), .S1(n1486), 
        .Y(n1280) );
  MXI4X1 U2285 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n2018), .S1(n1987), .Y(
        n1673) );
  MXI4X1 U2286 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n2018), .S1(n1987), .Y(
        n1677) );
  MXI4X1 U2287 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n2018), .S1(n1987), 
        .Y(n1681) );
  MXI4X1 U2288 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n2019), .S1(n1987), 
        .Y(n1685) );
  MXI4X1 U2289 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1689) );
  MXI4X1 U2290 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n2019), .S1(n1987), 
        .Y(n1693) );
  MXI4X1 U2291 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1697) );
  MXI4X1 U2292 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n2019), .S1(n1987), 
        .Y(n1701) );
  MXI4X1 U2293 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n2020), .S1(n1986), 
        .Y(n1705) );
  MXI4X1 U2294 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n2020), .S1(n1986), 
        .Y(n1709) );
  MXI4X1 U2295 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1717) );
  MXI4X1 U2296 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n2020), .S1(n1986), 
        .Y(n1713) );
  MXI4X1 U2297 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n2021), .S1(n1986), 
        .Y(n1725) );
  MXI4X1 U2298 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n2020), .S1(n1986), 
        .Y(n1721) );
  MXI4X1 U2299 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n2008), .S1(n1982), 
        .Y(n1733) );
  MXI4X1 U2300 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n2008), .S1(n1981), 
        .Y(n1729) );
  MXI4X1 U2301 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1741) );
  MXI4X1 U2302 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n2008), .S1(n1982), 
        .Y(n1737) );
  MXI4X1 U2303 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n2009), .S1(n1982), 
        .Y(n1749) );
  MXI4X1 U2304 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n2008), .S1(n1982), 
        .Y(n1745) );
  MXI4X1 U2305 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1757) );
  MXI4X1 U2306 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n2009), .S1(n1982), 
        .Y(n1753) );
  MXI4X1 U2307 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1765) );
  MXI4X1 U2308 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n2009), .S1(n1982), 
        .Y(n1761) );
  MXI4X1 U2309 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n2010), .S1(n1983), 
        .Y(n1773) );
  MXI4X1 U2310 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n2010), .S1(n1982), 
        .Y(n1769) );
  MXI4X1 U2311 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1781) );
  MXI4X1 U2312 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n2010), .S1(n1983), 
        .Y(n1777) );
  MXI4X1 U2313 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n2011), .S1(n1983), 
        .Y(n1789) );
  MXI4X1 U2314 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n2010), .S1(n1983), 
        .Y(n1785) );
  MXI4X1 U2315 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1797) );
  MXI4X1 U2316 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n2011), .S1(n1983), 
        .Y(n1793) );
  MXI4X1 U2317 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n2012), .S1(n1983), 
        .Y(n1805) );
  MXI4X1 U2318 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n2011), .S1(n1983), 
        .Y(n1801) );
  MXI4X1 U2319 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1813) );
  MXI4X1 U2320 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n2012), .S1(n1983), 
        .Y(n1809) );
  MXI4X1 U2321 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1821) );
  MXI4X1 U2322 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n2012), .S1(n1984), 
        .Y(n1817) );
  MXI4X1 U2323 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1829) );
  MXI4X1 U2324 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n2013), .S1(n1984), 
        .Y(n1825) );
  MXI4X1 U2325 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1837) );
  MXI4X1 U2326 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n2013), .S1(n1984), 
        .Y(n1833) );
  MXI4X1 U2327 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n2014), .S1(n1984), 
        .Y(n1845) );
  MXI4X1 U2328 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n2013), .S1(n1984), 
        .Y(n1841) );
  MXI4X1 U2329 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n2011), .S1(n1983), 
        .Y(n1853) );
  MXI4X1 U2330 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n2014), .S1(n1984), 
        .Y(n1849) );
  MX4X1 U2331 ( .A(n1298), .B(n1296), .C(n1297), .D(n1295), .S0(n1464), .S1(
        n1472), .Y(n1088) );
  MX4X1 U2332 ( .A(n1302), .B(n1300), .C(n1301), .D(n1299), .S0(n1464), .S1(
        n1472), .Y(n1087) );
  MXI4X1 U2333 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1295) );
  MX4X1 U2334 ( .A(n1306), .B(n1304), .C(n1305), .D(n1303), .S0(n1464), .S1(
        n1472), .Y(n1090) );
  MX4X1 U2335 ( .A(n1310), .B(n1308), .C(n1309), .D(n1307), .S0(n1464), .S1(
        n1473), .Y(n1089) );
  MXI4X1 U2336 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1514), .S1(n1486), 
        .Y(n1303) );
  MX4X1 U2337 ( .A(n1346), .B(n1344), .C(n1345), .D(n1343), .S0(n1465), .S1(
        n1473), .Y(n1100) );
  MX4X1 U2338 ( .A(n1350), .B(n1348), .C(n1349), .D(n1347), .S0(n1465), .S1(
        n1473), .Y(n1099) );
  MXI4X1 U2339 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1516), .S1(n1487), 
        .Y(n1343) );
  MXI2X1 U2340 ( .A(n1091), .B(n1092), .S0(n1457), .Y(ReadData1[26]) );
  MX4X1 U2341 ( .A(n1314), .B(n1312), .C(n1313), .D(n1311), .S0(n1465), .S1(
        n1473), .Y(n1092) );
  MX4X1 U2342 ( .A(n1318), .B(n1316), .C(n1317), .D(n1315), .S0(n1465), .S1(
        n1473), .Y(n1091) );
  MXI4X1 U2343 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1311) );
  MXI2X1 U2344 ( .A(n1093), .B(n1094), .S0(n1457), .Y(ReadData1[27]) );
  MX4X1 U2345 ( .A(n1322), .B(n1320), .C(n1321), .D(n1319), .S0(n1465), .S1(
        n1473), .Y(n1094) );
  MX4X1 U2346 ( .A(n1326), .B(n1324), .C(n1325), .D(n1323), .S0(n1465), .S1(
        n1473), .Y(n1093) );
  MXI4X1 U2347 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1319) );
  MXI2X1 U2348 ( .A(n1097), .B(n1098), .S0(n1457), .Y(ReadData1[29]) );
  MX4X1 U2349 ( .A(n1338), .B(n1336), .C(n1337), .D(n1335), .S0(n1465), .S1(
        n1473), .Y(n1098) );
  MX4X1 U2350 ( .A(n1342), .B(n1340), .C(n1341), .D(n1339), .S0(n1465), .S1(
        n1473), .Y(n1097) );
  MXI4X1 U2351 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1335) );
  MXI2X1 U2352 ( .A(n1095), .B(n1096), .S0(n1457), .Y(ReadData1[28]) );
  MX4X1 U2353 ( .A(n1330), .B(n1328), .C(n1329), .D(n1327), .S0(n1465), .S1(
        n1473), .Y(n1096) );
  MX4X1 U2354 ( .A(n1334), .B(n1332), .C(n1333), .D(n1331), .S0(n1465), .S1(
        n1473), .Y(n1095) );
  MXI4X1 U2355 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1327) );
  MXI2X1 U2356 ( .A(n1101), .B(n1102), .S0(n1457), .Y(ReadData1[31]) );
  MX4X1 U2357 ( .A(n1354), .B(n1352), .C(n1353), .D(n1351), .S0(n1465), .S1(
        n1473), .Y(n1102) );
  MX4X1 U2358 ( .A(n1358), .B(n1356), .C(n1357), .D(n1355), .S0(n1465), .S1(
        n1473), .Y(n1101) );
  MXI4X1 U2359 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1517), .S1(n1487), 
        .Y(n1351) );
  MXI2X1 U2360 ( .A(n1085), .B(n1086), .S0(n1457), .Y(ReadData1[23]) );
  MX4X1 U2361 ( .A(n1290), .B(n1288), .C(n1289), .D(n1287), .S0(n1464), .S1(
        n1472), .Y(n1086) );
  MX4X1 U2362 ( .A(n1294), .B(n1292), .C(n1293), .D(n1291), .S0(n1464), .S1(
        n1472), .Y(n1085) );
  MXI4X1 U2363 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1513), .S1(n1486), 
        .Y(n1287) );
  NAND2BX1 U2364 ( .AN(n1385), .B(n1384), .Y(n1294) );
  MXI2X1 U2365 ( .A(n2388), .B(n1383), .S0(n1527), .Y(n1384) );
  OAI22XL U2366 ( .A0(n1495), .A1(n1525), .B0(n1493), .B1(\register[1][23] ), 
        .Y(n1385) );
  NOR2BX1 U2367 ( .AN(n1491), .B(\register[3][23] ), .Y(n1383) );
  NAND2BX1 U2368 ( .AN(n1379), .B(n1378), .Y(n1310) );
  MXI2X1 U2369 ( .A(n2390), .B(n1377), .S0(n1527), .Y(n1378) );
  OAI22XL U2370 ( .A0(n1495), .A1(n1525), .B0(n1494), .B1(\register[1][25] ), 
        .Y(n1379) );
  NOR2BX1 U2371 ( .AN(n1491), .B(\register[3][25] ), .Y(n1377) );
  NAND2BX1 U2372 ( .AN(n1376), .B(n1375), .Y(n1318) );
  MXI2X1 U2373 ( .A(n2391), .B(n1374), .S0(n1527), .Y(n1375) );
  OAI22XL U2374 ( .A0(n1495), .A1(n1526), .B0(n1493), .B1(\register[1][26] ), 
        .Y(n1376) );
  NOR2BX1 U2375 ( .AN(n1491), .B(\register[3][26] ), .Y(n1374) );
  NAND2BX1 U2376 ( .AN(n1373), .B(n1372), .Y(n1326) );
  MXI2X1 U2377 ( .A(n2392), .B(n1371), .S0(n1527), .Y(n1372) );
  OAI22XL U2378 ( .A0(n1496), .A1(n1526), .B0(n1494), .B1(\register[1][27] ), 
        .Y(n1373) );
  NOR2BX1 U2379 ( .AN(n1491), .B(\register[3][27] ), .Y(n1371) );
  NAND2BX1 U2380 ( .AN(n1364), .B(n1363), .Y(n1350) );
  MXI2X1 U2381 ( .A(n2395), .B(n1362), .S0(n1528), .Y(n1363) );
  OAI22XL U2382 ( .A0(n1496), .A1(n1526), .B0(n1493), .B1(\register[1][30] ), 
        .Y(n1364) );
  NOR2BX1 U2383 ( .AN(n1491), .B(\register[3][30] ), .Y(n1362) );
  NAND2BX1 U2384 ( .AN(n1370), .B(n1369), .Y(n1334) );
  MXI2X1 U2385 ( .A(n2393), .B(n1368), .S0(n1528), .Y(n1369) );
  OAI22XL U2386 ( .A0(n1496), .A1(n1525), .B0(n1494), .B1(\register[1][28] ), 
        .Y(n1370) );
  NOR2BX1 U2387 ( .AN(n1491), .B(\register[3][28] ), .Y(n1368) );
  NAND2BX1 U2388 ( .AN(n1367), .B(n1366), .Y(n1342) );
  MXI2X1 U2389 ( .A(n2394), .B(n1365), .S0(n1528), .Y(n1366) );
  OAI22XL U2390 ( .A0(n1496), .A1(n1526), .B0(n1494), .B1(\register[1][29] ), 
        .Y(n1367) );
  NOR2BX1 U2391 ( .AN(n1491), .B(\register[3][29] ), .Y(n1365) );
  NAND2BX1 U2392 ( .AN(n1361), .B(n1360), .Y(n1358) );
  MXI2X1 U2393 ( .A(n2396), .B(n1359), .S0(n1528), .Y(n1360) );
  OAI22XL U2394 ( .A0(n1496), .A1(n1525), .B0(n1494), .B1(\register[1][31] ), 
        .Y(n1361) );
  NOR2BX1 U2395 ( .AN(n1491), .B(\register[3][31] ), .Y(n1359) );
  NAND2BX1 U2396 ( .AN(n1382), .B(n1381), .Y(n1302) );
  MXI2X1 U2397 ( .A(n2389), .B(n1380), .S0(n1526), .Y(n1381) );
  OAI22XL U2398 ( .A0(n1496), .A1(n1526), .B0(n1493), .B1(\register[1][24] ), 
        .Y(n1382) );
  NOR2BX1 U2399 ( .AN(n1491), .B(\register[3][24] ), .Y(n1380) );
  MXI4X1 U2400 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1514), .S1(n1486), .Y(
        n1293) );
  MXI4X1 U2401 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1514), .S1(n1486), 
        .Y(n1289) );
  MXI4X1 U2402 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1514), .S1(n1486), .Y(
        n1301) );
  MXI4X1 U2403 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1297) );
  MXI4X1 U2404 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1515), .S1(n1486), .Y(
        n1309) );
  MXI4X1 U2405 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1514), .S1(n1486), 
        .Y(n1305) );
  MXI4X1 U2406 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1515), .S1(n1487), .Y(
        n1317) );
  MXI4X1 U2407 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1313) );
  MXI4X1 U2408 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1515), .S1(n1487), .Y(
        n1325) );
  MXI4X1 U2409 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1321) );
  MXI4X1 U2410 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1517), .S1(n1487), .Y(
        n1349) );
  MXI4X1 U2411 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1516), .S1(n1487), 
        .Y(n1345) );
  MXI4X1 U2412 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1516), .S1(n1487), .Y(
        n1333) );
  MXI4X1 U2413 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1329) );
  MXI4X1 U2414 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1516), .S1(n1487), .Y(
        n1341) );
  MXI4X1 U2415 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1337) );
  MXI4X1 U2416 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1524), .S1(n1489), .Y(
        n1357) );
  MXI4X1 U2417 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1517), .S1(n1487), 
        .Y(n1353) );
  MXI4X1 U2418 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1514), .S1(n1486), 
        .Y(n1290) );
  MXI4X1 U2419 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1298) );
  MXI4X1 U2420 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1514), .S1(n1486), 
        .Y(n1306) );
  MXI4X1 U2421 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1314) );
  MXI4X1 U2422 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1322) );
  MXI4X1 U2423 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1517), .S1(n1487), 
        .Y(n1346) );
  MXI4X1 U2424 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1330) );
  MXI4X1 U2425 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1338) );
  MXI4X1 U2426 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1517), .S1(n1487), 
        .Y(n1354) );
  MXI4X1 U2427 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1514), .S1(n1486), 
        .Y(n1291) );
  MXI4X1 U2428 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1299) );
  MXI4X1 U2429 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1515), .S1(n1486), 
        .Y(n1307) );
  MXI4X1 U2430 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1315) );
  MXI4X1 U2431 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1323) );
  MXI4X1 U2432 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1517), .S1(n1487), 
        .Y(n1347) );
  MXI4X1 U2433 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1331) );
  MXI4X1 U2434 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1339) );
  MXI4X1 U2435 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1517), .S1(n1487), 
        .Y(n1355) );
  MXI4X1 U2436 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1514), .S1(n1486), 
        .Y(n1292) );
  MXI4X1 U2437 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1513), .S1(n1486), 
        .Y(n1288) );
  MXI4X1 U2438 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1300) );
  MXI4X1 U2439 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1514), .S1(n1486), 
        .Y(n1296) );
  MXI4X1 U2440 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1515), .S1(n1486), 
        .Y(n1308) );
  MXI4X1 U2441 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1514), .S1(n1486), 
        .Y(n1304) );
  MXI4X1 U2442 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1316) );
  MXI4X1 U2443 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1515), .S1(n1486), 
        .Y(n1312) );
  MXI4X1 U2444 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1324) );
  MXI4X1 U2445 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1515), .S1(n1487), 
        .Y(n1320) );
  MXI4X1 U2446 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1517), .S1(n1487), 
        .Y(n1348) );
  MXI4X1 U2447 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1516), .S1(n1487), 
        .Y(n1344) );
  MXI4X1 U2448 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1332) );
  MXI4X1 U2449 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1516), .S1(n1487), 
        .Y(n1328) );
  MXI4X1 U2450 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1340) );
  MXI4X1 U2451 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1516), .S1(n1487), 
        .Y(n1336) );
  MXI4X1 U2452 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1514), .S1(n1486), 
        .Y(n1356) );
  MXI4X1 U2453 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1517), .S1(n1487), 
        .Y(n1352) );
  NOR2BX1 U2454 ( .AN(RegWrite), .B(n2350), .Y(n53) );
  CLKBUFX3 U2455 ( .A(n1458), .Y(n1455) );
  CLKBUFX3 U2456 ( .A(N17), .Y(n1458) );
  CLKBUFX3 U2457 ( .A(n1955), .Y(n1952) );
  CLKBUFX3 U2458 ( .A(N22), .Y(n1955) );
  CLKBUFX3 U2459 ( .A(n1474), .Y(n1469) );
  CLKBUFX3 U2460 ( .A(N15), .Y(n1474) );
  CLKBUFX3 U2461 ( .A(N17), .Y(n1459) );
  CLKBUFX3 U2462 ( .A(N15), .Y(n1475) );
  CLKBUFX3 U2463 ( .A(N15), .Y(n1476) );
  CLKBUFX3 U2464 ( .A(N22), .Y(n1956) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  XOR3X1 U2_31 ( .A(A[31]), .B(n9), .C(carry[31]), .Y(DIFF[31]) );
  ADDFXL U2_30 ( .A(A[30]), .B(n10), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n12), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n13), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n14), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n15), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n16), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n17), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n18), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n19), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n20), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n21), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n23), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n24), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n25), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n26), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n27), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n28), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n29), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n30), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n31), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n32), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n2), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n3), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n4), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n5), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n6), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n8), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n22), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  INVXL U1 ( .A(B[15]), .Y(n27) );
  INVXL U2 ( .A(B[6]), .Y(n5) );
  INVXL U3 ( .A(B[7]), .Y(n4) );
  INVXL U4 ( .A(B[14]), .Y(n28) );
  NAND2BX1 U5 ( .AN(n33), .B(n1), .Y(carry[1]) );
  INVXL U6 ( .A(B[8]), .Y(n3) );
  INVXL U7 ( .A(B[9]), .Y(n2) );
  INVXL U8 ( .A(B[10]), .Y(n32) );
  INVXL U9 ( .A(B[11]), .Y(n31) );
  INVXL U10 ( .A(B[12]), .Y(n30) );
  INVXL U11 ( .A(B[13]), .Y(n29) );
  INVXL U12 ( .A(B[16]), .Y(n26) );
  INVXL U13 ( .A(B[0]), .Y(n33) );
  XNOR2X1 U14 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U15 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U16 ( .A(B[1]), .Y(n22) );
  CLKINVX1 U17 ( .A(B[2]), .Y(n11) );
  CLKINVX1 U18 ( .A(B[3]), .Y(n8) );
  CLKINVX1 U19 ( .A(B[4]), .Y(n7) );
  CLKINVX1 U20 ( .A(B[5]), .Y(n6) );
  CLKINVX1 U21 ( .A(B[17]), .Y(n25) );
  CLKINVX1 U22 ( .A(B[18]), .Y(n24) );
  CLKINVX1 U23 ( .A(B[19]), .Y(n23) );
  CLKINVX1 U24 ( .A(B[20]), .Y(n21) );
  CLKINVX1 U25 ( .A(B[21]), .Y(n20) );
  CLKINVX1 U26 ( .A(B[22]), .Y(n19) );
  CLKINVX1 U27 ( .A(B[23]), .Y(n18) );
  CLKINVX1 U28 ( .A(B[24]), .Y(n17) );
  CLKINVX1 U29 ( .A(B[25]), .Y(n16) );
  CLKINVX1 U30 ( .A(B[26]), .Y(n15) );
  CLKINVX1 U31 ( .A(B[27]), .Y(n14) );
  CLKINVX1 U32 ( .A(B[28]), .Y(n13) );
  CLKINVX1 U33 ( .A(B[29]), .Y(n12) );
  CLKINVX1 U34 ( .A(B[30]), .Y(n10) );
  CLKINVX1 U35 ( .A(B[31]), .Y(n9) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110;

  OAI221X1 U1 ( .A0(A[10]), .A1(n25), .B0(A[11]), .B1(n24), .C0(n96), .Y(n95)
         );
  AND4X4 U2 ( .A(n38), .B(n39), .C(n40), .D(n41), .Y(EQ) );
  NOR4BBX1 U3 ( .AN(n73), .BN(n74), .C(LT), .D(n75), .Y(n39) );
  OAI221X1 U4 ( .A0(A[28]), .A1(n12), .B0(A[29]), .B1(n11), .C0(n78), .Y(n77)
         );
  OAI211X1 U5 ( .A0(n79), .A1(n80), .B0(n49), .C0(n53), .Y(n78) );
  OAI221X1 U6 ( .A0(A[12]), .A1(n23), .B0(A[13]), .B1(n22), .C0(n94), .Y(n93)
         );
  OAI221X1 U7 ( .A0(A[20]), .A1(n17), .B0(A[21]), .B1(n16), .C0(n86), .Y(n85)
         );
  OAI211X1 U8 ( .A0(n87), .A1(n88), .B0(n58), .C0(n61), .Y(n86) );
  OR2X2 U9 ( .A(n2), .B(n3), .Y(LT) );
  AOI221XL U10 ( .A0(B[7]), .A1(n33), .B0(B[6]), .B1(n34), .C0(n101), .Y(n99)
         );
  AOI221XL U11 ( .A0(B[25]), .A1(n27), .B0(B[24]), .B1(n28), .C0(n82), .Y(n81)
         );
  AO21X2 U12 ( .A0(n37), .A1(n108), .B0(B[1]), .Y(n109) );
  AOI32X1 U13 ( .A0(n7), .A1(n74), .A2(n106), .B0(B[4]), .B1(n36), .Y(n102) );
  AOI32X1 U14 ( .A0(n66), .A1(n67), .A2(n93), .B0(B[14]), .B1(n32), .Y(n91) );
  AOI32X1 U15 ( .A0(n56), .A1(n57), .A2(n85), .B0(B[22]), .B1(n29), .Y(n83) );
  OAI221X1 U16 ( .A0(A[2]), .A1(n10), .B0(A[3]), .B1(n8), .C0(n107), .Y(n106)
         );
  NOR2BX1 U17 ( .AN(B[0]), .B(A[0]), .Y(n108) );
  OAI211XL U18 ( .A0(n97), .A1(n98), .B0(n70), .C0(n71), .Y(n96) );
  AOI32XL U19 ( .A0(n47), .A1(n48), .A2(n77), .B0(B[30]), .B1(n26), .Y(n76) );
  NOR2X1 U20 ( .A(n33), .B(B[7]), .Y(n100) );
  NAND4BXL U21 ( .AN(n65), .B(n66), .C(n67), .D(n68), .Y(n64) );
  NAND4XL U22 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n63) );
  INVX1 U23 ( .A(n72), .Y(n5) );
  OAI211XL U24 ( .A0(n108), .A1(n37), .B0(n109), .C0(n73), .Y(n107) );
  NOR2XL U25 ( .A(n35), .B(B[5]), .Y(n104) );
  NOR2BXL U26 ( .AN(A[15]), .B(B[15]), .Y(n65) );
  NAND2XL U27 ( .A(A[11]), .B(n24), .Y(n69) );
  NAND2XL U28 ( .A(A[13]), .B(n22), .Y(n67) );
  NAND2XL U29 ( .A(A[3]), .B(n8), .Y(n74) );
  INVX1 U30 ( .A(B[8]), .Y(n6) );
  INVX1 U31 ( .A(B[9]), .Y(n4) );
  INVX1 U32 ( .A(B[11]), .Y(n24) );
  INVX1 U33 ( .A(B[13]), .Y(n22) );
  INVX1 U34 ( .A(B[10]), .Y(n25) );
  INVX1 U35 ( .A(B[12]), .Y(n23) );
  NOR2BXL U36 ( .AN(A[0]), .B(B[0]), .Y(n50) );
  NOR2X1 U37 ( .A(A[31]), .B(n9), .Y(n2) );
  NOR2X1 U38 ( .A(n75), .B(n76), .Y(n3) );
  CLKINVX1 U39 ( .A(B[18]), .Y(n21) );
  CLKINVX1 U40 ( .A(B[19]), .Y(n19) );
  CLKINVX1 U41 ( .A(B[21]), .Y(n16) );
  CLKINVX1 U42 ( .A(B[20]), .Y(n17) );
  CLKINVX1 U43 ( .A(n62), .Y(n20) );
  CLKINVX1 U44 ( .A(B[26]), .Y(n15) );
  CLKINVX1 U45 ( .A(B[27]), .Y(n13) );
  CLKINVX1 U46 ( .A(B[29]), .Y(n11) );
  CLKINVX1 U47 ( .A(B[28]), .Y(n12) );
  CLKINVX1 U48 ( .A(B[31]), .Y(n9) );
  CLKINVX1 U49 ( .A(n54), .Y(n14) );
  CLKINVX1 U50 ( .A(n110), .Y(n7) );
  CLKINVX1 U51 ( .A(A[4]), .Y(n36) );
  CLKINVX1 U52 ( .A(A[5]), .Y(n35) );
  CLKINVX1 U53 ( .A(A[1]), .Y(n37) );
  CLKINVX1 U54 ( .A(A[7]), .Y(n33) );
  CLKINVX1 U55 ( .A(A[6]), .Y(n34) );
  CLKINVX1 U56 ( .A(B[3]), .Y(n8) );
  CLKINVX1 U57 ( .A(B[2]), .Y(n10) );
  CLKINVX1 U58 ( .A(A[17]), .Y(n30) );
  CLKINVX1 U59 ( .A(A[16]), .Y(n31) );
  CLKINVX1 U60 ( .A(A[14]), .Y(n32) );
  CLKINVX1 U61 ( .A(A[22]), .Y(n29) );
  CLKINVX1 U62 ( .A(B[1]), .Y(n18) );
  CLKINVX1 U63 ( .A(A[25]), .Y(n27) );
  CLKINVX1 U64 ( .A(A[24]), .Y(n28) );
  CLKINVX1 U65 ( .A(A[30]), .Y(n26) );
  NOR4X1 U66 ( .A(n42), .B(n43), .C(n44), .D(n45), .Y(n41) );
  NAND4X1 U67 ( .A(n46), .B(n47), .C(n48), .D(n49), .Y(n45) );
  OAI22XL U68 ( .A0(A[1]), .A1(n50), .B0(n50), .B1(n18), .Y(n46) );
  NAND4BBXL U69 ( .AN(n51), .BN(n52), .C(n53), .D(n54), .Y(n44) );
  NAND4BX1 U70 ( .AN(n55), .B(n56), .C(n57), .D(n58), .Y(n43) );
  NAND4BBXL U71 ( .AN(n59), .BN(n60), .C(n61), .D(n62), .Y(n42) );
  NOR2X1 U72 ( .A(n63), .B(n64), .Y(n40) );
  NAND2X1 U73 ( .A(A[27]), .B(n13), .Y(n53) );
  NAND2X1 U74 ( .A(A[28]), .B(n12), .Y(n49) );
  OAI32X1 U75 ( .A0(n81), .A1(n51), .A2(n14), .B0(A[26]), .B1(n15), .Y(n80) );
  NAND2X1 U76 ( .A(A[26]), .B(n15), .Y(n54) );
  NOR2X1 U77 ( .A(n27), .B(B[25]), .Y(n51) );
  AOI211X1 U78 ( .A0(n83), .A1(n84), .B0(n55), .C0(n52), .Y(n82) );
  NOR2X1 U79 ( .A(n28), .B(B[24]), .Y(n52) );
  NOR2BX1 U80 ( .AN(A[23]), .B(B[23]), .Y(n55) );
  NAND2BX1 U81 ( .AN(A[23]), .B(B[23]), .Y(n84) );
  NAND2X1 U82 ( .A(A[19]), .B(n19), .Y(n61) );
  NAND2X1 U83 ( .A(A[20]), .B(n17), .Y(n58) );
  OAI32X1 U84 ( .A0(n89), .A1(n59), .A2(n20), .B0(A[18]), .B1(n21), .Y(n88) );
  NAND2X1 U85 ( .A(A[18]), .B(n21), .Y(n62) );
  NOR2X1 U86 ( .A(n30), .B(B[17]), .Y(n59) );
  AOI221XL U87 ( .A0(B[17]), .A1(n30), .B0(B[16]), .B1(n31), .C0(n90), .Y(n89)
         );
  AOI211X1 U88 ( .A0(n91), .A1(n92), .B0(n65), .C0(n60), .Y(n90) );
  NOR2X1 U89 ( .A(n31), .B(B[16]), .Y(n60) );
  NAND2BX1 U90 ( .AN(A[15]), .B(B[15]), .Y(n92) );
  NAND3X1 U91 ( .A(n68), .B(n69), .C(n95), .Y(n94) );
  NAND2X1 U92 ( .A(A[9]), .B(n4), .Y(n71) );
  NAND2X1 U93 ( .A(A[10]), .B(n25), .Y(n70) );
  OAI32X1 U94 ( .A0(n99), .A1(n100), .A2(n5), .B0(A[8]), .B1(n6), .Y(n98) );
  NAND2X1 U95 ( .A(A[8]), .B(n6), .Y(n72) );
  AOI211X1 U96 ( .A0(n102), .A1(n103), .B0(n104), .C0(n105), .Y(n101) );
  NAND2X1 U97 ( .A(B[5]), .B(n35), .Y(n103) );
  NOR2X1 U98 ( .A(A[9]), .B(n4), .Y(n97) );
  NAND2X1 U99 ( .A(A[12]), .B(n23), .Y(n68) );
  OR2X1 U100 ( .A(B[14]), .B(n32), .Y(n66) );
  NOR2X1 U101 ( .A(A[19]), .B(n19), .Y(n87) );
  NAND2X1 U102 ( .A(A[21]), .B(n16), .Y(n57) );
  OR2X1 U103 ( .A(B[22]), .B(n29), .Y(n56) );
  NOR2X1 U104 ( .A(A[27]), .B(n13), .Y(n79) );
  OR2X1 U105 ( .A(B[30]), .B(n26), .Y(n48) );
  NAND2X1 U106 ( .A(A[29]), .B(n11), .Y(n47) );
  NOR2BX1 U107 ( .AN(A[31]), .B(B[31]), .Y(n75) );
  NAND2X1 U108 ( .A(A[2]), .B(n10), .Y(n73) );
  NOR4X1 U109 ( .A(n110), .B(n104), .C(n105), .D(n100), .Y(n38) );
  NOR2X1 U110 ( .A(n34), .B(B[6]), .Y(n105) );
  NOR2X1 U111 ( .A(n36), .B(B[4]), .Y(n110) );
endmodule


module alu ( ctrl, x, y, zero, out );
  input [3:0] ctrl;
  input [31:0] x;
  input [31:0] y;
  output [31:0] out;
  output zero;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N134, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n185, n186, n187, n188;

  alu_DW01_sub_0 sub_248 ( .A(x), .B(y), .CI(1'b0), .DIFF({N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70}) );
  alu_DW01_add_0 add_246 ( .A(x), .B(y), .CI(1'b0), .SUM({N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38})
         );
  alu_DW01_cmp6_0 r302 ( .A(x), .B(y), .TC(1'b0), .LT(N134), .EQ(N200) );
  TLATX1 \prev_out_reg[31]  ( .G(N167), .D(N199), .Q(out[31]) );
  TLATX1 \prev_out_reg[30]  ( .G(N167), .D(N198), .Q(out[30]) );
  TLATX1 \prev_out_reg[29]  ( .G(N167), .D(N197), .Q(out[29]) );
  TLATX1 \prev_out_reg[28]  ( .G(N167), .D(N196), .Q(out[28]) );
  TLATX1 \prev_out_reg[27]  ( .G(N167), .D(N195), .Q(out[27]) );
  TLATX1 \prev_out_reg[26]  ( .G(N167), .D(N194), .Q(out[26]) );
  TLATX1 \prev_out_reg[25]  ( .G(N167), .D(N193), .Q(out[25]) );
  TLATX1 \prev_out_reg[24]  ( .G(N167), .D(N192), .Q(out[24]) );
  TLATX1 \prev_out_reg[23]  ( .G(N167), .D(N191), .Q(out[23]) );
  TLATX1 \prev_out_reg[22]  ( .G(N167), .D(N190), .Q(out[22]) );
  TLATX1 \prev_out_reg[21]  ( .G(N167), .D(N189), .Q(out[21]) );
  TLATX1 \prev_out_reg[20]  ( .G(N167), .D(N188), .Q(out[20]) );
  TLATX1 \prev_out_reg[19]  ( .G(N167), .D(N187), .Q(out[19]) );
  TLATX1 \prev_out_reg[18]  ( .G(N167), .D(N186), .Q(out[18]) );
  TLATX1 \prev_out_reg[17]  ( .G(N167), .D(N185), .Q(out[17]) );
  TLATX1 \prev_out_reg[16]  ( .G(N167), .D(N184), .Q(out[16]) );
  TLATX1 \prev_out_reg[15]  ( .G(N167), .D(N183), .Q(out[15]) );
  TLATX1 \prev_out_reg[14]  ( .G(N167), .D(N182), .Q(out[14]) );
  TLATX1 \prev_out_reg[13]  ( .G(N167), .D(N181), .Q(out[13]) );
  TLATX1 \prev_out_reg[12]  ( .G(N167), .D(N180), .Q(out[12]) );
  TLATX1 \prev_out_reg[11]  ( .G(N167), .D(N179), .Q(out[11]) );
  TLATX1 \prev_out_reg[10]  ( .G(N167), .D(N178), .Q(out[10]) );
  TLATX1 \prev_out_reg[9]  ( .G(N167), .D(N177), .Q(out[9]) );
  TLATX1 \prev_out_reg[8]  ( .G(N167), .D(N176), .Q(out[8]) );
  TLATX1 \prev_out_reg[7]  ( .G(N167), .D(N175), .Q(out[7]) );
  TLATX1 \prev_out_reg[6]  ( .G(N167), .D(N174), .Q(out[6]) );
  TLATX1 \prev_out_reg[5]  ( .G(N167), .D(N173), .Q(out[5]) );
  TLATX1 \prev_out_reg[4]  ( .G(N167), .D(N172), .Q(out[4]) );
  TLATX1 \prev_out_reg[3]  ( .G(N167), .D(N171), .Q(out[3]) );
  TLATX1 \prev_out_reg[2]  ( .G(N167), .D(N170), .Q(out[2]) );
  TLATX1 \prev_out_reg[1]  ( .G(N167), .D(N169), .Q(out[1]) );
  TLATX1 \prev_out_reg[0]  ( .G(N167), .D(N168), .Q(out[0]) );
  TLATX1 prev_zero_reg ( .G(1'b1), .D(N200), .Q(zero) );
  AOI32XL U2 ( .A0(n187), .A1(n40), .A2(n85), .B0(y[1]), .B1(n177), .Y(n175)
         );
  AOI32XL U3 ( .A0(n69), .A1(n45), .A2(n4), .B0(y[15]), .B1(n135), .Y(n133) );
  INVXL U7 ( .A(y[15]), .Y(n45) );
  INVXL U8 ( .A(y[16]), .Y(n44) );
  CLKINVX1 U9 ( .A(n14), .Y(n15) );
  AOI32XL U10 ( .A0(n76), .A1(n21), .A2(n85), .B0(y[8]), .B1(n156), .Y(n154)
         );
  INVXL U11 ( .A(y[8]), .Y(n21) );
  AOI32XL U12 ( .A0(n75), .A1(n20), .A2(n4), .B0(y[9]), .B1(n153), .Y(n151) );
  INVXL U13 ( .A(y[9]), .Y(n20) );
  AOI32XL U14 ( .A0(n74), .A1(n50), .A2(n85), .B0(y[10]), .B1(n150), .Y(n148)
         );
  INVXL U15 ( .A(y[10]), .Y(n50) );
  AOI32XL U16 ( .A0(n73), .A1(n49), .A2(n4), .B0(y[11]), .B1(n147), .Y(n145)
         );
  INVXL U17 ( .A(y[11]), .Y(n49) );
  AOI32XL U18 ( .A0(n72), .A1(n48), .A2(n85), .B0(y[12]), .B1(n144), .Y(n142)
         );
  INVXL U19 ( .A(y[12]), .Y(n48) );
  AOI32XL U20 ( .A0(n71), .A1(n47), .A2(n4), .B0(y[13]), .B1(n141), .Y(n139)
         );
  INVXL U21 ( .A(y[13]), .Y(n47) );
  AOI32XL U22 ( .A0(n70), .A1(n46), .A2(n85), .B0(y[14]), .B1(n138), .Y(n136)
         );
  INVXL U23 ( .A(y[14]), .Y(n46) );
  AOI32XL U24 ( .A0(n78), .A1(n23), .A2(n85), .B0(y[6]), .B1(n162), .Y(n160)
         );
  INVXL U25 ( .A(y[6]), .Y(n23) );
  AOI32XL U26 ( .A0(n77), .A1(n22), .A2(n4), .B0(y[7]), .B1(n159), .Y(n157) );
  INVXL U27 ( .A(y[7]), .Y(n22) );
  INVXL U28 ( .A(x[8]), .Y(n76) );
  INVXL U29 ( .A(x[9]), .Y(n75) );
  INVXL U30 ( .A(x[3]), .Y(n185) );
  INVXL U31 ( .A(x[11]), .Y(n73) );
  INVXL U32 ( .A(x[13]), .Y(n71) );
  INVXL U33 ( .A(x[2]), .Y(n186) );
  INVXL U34 ( .A(x[10]), .Y(n74) );
  INVXL U35 ( .A(x[12]), .Y(n72) );
  INVXL U36 ( .A(x[15]), .Y(n69) );
  NOR4X1 U37 ( .A(n18), .B(n19), .C(ctrl[0]), .D(ctrl[3]), .Y(n84) );
  INVXL U38 ( .A(y[0]), .Y(n51) );
  AOI33XL U39 ( .A0(N134), .A1(ctrl[1]), .A2(n182), .B0(n188), .B1(n51), .B2(
        n85), .Y(n179) );
  CLKBUFX3 U40 ( .A(n16), .Y(n6) );
  CLKBUFX3 U41 ( .A(n16), .Y(n5) );
  CLKBUFX3 U42 ( .A(n16), .Y(n7) );
  CLKINVX1 U43 ( .A(n181), .Y(n16) );
  OAI21XL U44 ( .A0(n8), .A1(n187), .B0(n81), .Y(n177) );
  OAI21XL U45 ( .A0(n8), .A1(n80), .B0(n14), .Y(n168) );
  OAI21XL U46 ( .A0(n8), .A1(n79), .B0(n81), .Y(n165) );
  OAI21XL U47 ( .A0(n8), .A1(n78), .B0(n14), .Y(n162) );
  OAI21XL U48 ( .A0(n9), .A1(n77), .B0(n81), .Y(n159) );
  OAI21XL U49 ( .A0(n9), .A1(n70), .B0(n81), .Y(n138) );
  OAI21XL U50 ( .A0(n9), .A1(n68), .B0(n14), .Y(n132) );
  OAI21XL U51 ( .A0(n9), .A1(n67), .B0(n14), .Y(n129) );
  OAI21XL U52 ( .A0(n9), .A1(n62), .B0(n14), .Y(n114) );
  OAI21XL U53 ( .A0(n9), .A1(n60), .B0(n81), .Y(n108) );
  OAI21XL U54 ( .A0(n10), .A1(n59), .B0(n81), .Y(n105) );
  OAI21XL U55 ( .A0(n10), .A1(n54), .B0(n14), .Y(n90) );
  OAI21XL U56 ( .A0(n8), .A1(n76), .B0(n14), .Y(n156) );
  OAI21XL U57 ( .A0(n8), .A1(n75), .B0(n81), .Y(n153) );
  OAI21XL U58 ( .A0(n9), .A1(n66), .B0(n81), .Y(n126) );
  OAI21XL U59 ( .A0(n10), .A1(n58), .B0(n14), .Y(n102) );
  OAI21XL U60 ( .A0(n8), .A1(n186), .B0(n14), .Y(n174) );
  OAI21XL U61 ( .A0(n8), .A1(n185), .B0(n81), .Y(n171) );
  OAI21XL U62 ( .A0(n8), .A1(n74), .B0(n81), .Y(n150) );
  OAI21XL U63 ( .A0(n8), .A1(n73), .B0(n14), .Y(n147) );
  OAI21XL U64 ( .A0(n8), .A1(n72), .B0(n81), .Y(n144) );
  OAI21XL U65 ( .A0(n9), .A1(n71), .B0(n14), .Y(n141) );
  OAI21XL U66 ( .A0(n9), .A1(n65), .B0(n14), .Y(n123) );
  OAI21XL U67 ( .A0(n9), .A1(n64), .B0(n81), .Y(n120) );
  OAI21XL U68 ( .A0(n9), .A1(n63), .B0(n14), .Y(n117) );
  OAI21XL U69 ( .A0(n10), .A1(n57), .B0(n14), .Y(n99) );
  OAI21XL U70 ( .A0(n10), .A1(n56), .B0(n81), .Y(n96) );
  OAI21XL U71 ( .A0(n10), .A1(n55), .B0(n81), .Y(n93) );
  OAI21XL U72 ( .A0(n8), .A1(n53), .B0(n14), .Y(n86) );
  OAI21XL U73 ( .A0(n9), .A1(n69), .B0(n14), .Y(n135) );
  OAI21XL U74 ( .A0(n9), .A1(n61), .B0(n81), .Y(n111) );
  CLKBUFX3 U75 ( .A(n87), .Y(n8) );
  CLKBUFX3 U76 ( .A(n87), .Y(n9) );
  AOI2BB1X1 U77 ( .A0N(n10), .A1N(n188), .B0(n15), .Y(n178) );
  CLKBUFX3 U78 ( .A(n87), .Y(n10) );
  OAI211X1 U79 ( .A0(n53), .A1(n81), .B0(n82), .C0(n83), .Y(N199) );
  AOI32X1 U80 ( .A0(n53), .A1(n27), .A2(n4), .B0(y[31]), .B1(n86), .Y(n82) );
  AOI22X1 U81 ( .A0(N101), .A1(n11), .B0(N69), .B1(n5), .Y(n83) );
  CLKINVX1 U82 ( .A(y[31]), .Y(n27) );
  OAI211X1 U83 ( .A0(n14), .A1(n69), .B0(n133), .C0(n134), .Y(N183) );
  AOI22X1 U84 ( .A0(N85), .A1(n12), .B0(N53), .B1(n6), .Y(n134) );
  OAI211X1 U85 ( .A0(n81), .A1(n68), .B0(n130), .C0(n131), .Y(N184) );
  AOI32XL U86 ( .A0(n68), .A1(n44), .A2(n85), .B0(y[16]), .B1(n132), .Y(n130)
         );
  AOI22X1 U87 ( .A0(N86), .A1(n12), .B0(N54), .B1(n6), .Y(n131) );
  OAI211X1 U88 ( .A0(n14), .A1(n67), .B0(n127), .C0(n128), .Y(N185) );
  AOI32X1 U89 ( .A0(n67), .A1(n43), .A2(n4), .B0(y[17]), .B1(n129), .Y(n127)
         );
  AOI22X1 U90 ( .A0(N87), .A1(n12), .B0(N55), .B1(n6), .Y(n128) );
  CLKINVX1 U91 ( .A(y[17]), .Y(n43) );
  OAI211X1 U92 ( .A0(n81), .A1(n66), .B0(n124), .C0(n125), .Y(N186) );
  AOI32XL U93 ( .A0(n66), .A1(n42), .A2(n85), .B0(y[18]), .B1(n126), .Y(n124)
         );
  AOI22X1 U94 ( .A0(N88), .A1(n12), .B0(N56), .B1(n6), .Y(n125) );
  CLKINVX1 U95 ( .A(y[18]), .Y(n42) );
  OAI211X1 U96 ( .A0(n14), .A1(n65), .B0(n121), .C0(n122), .Y(N187) );
  AOI32X1 U97 ( .A0(n65), .A1(n41), .A2(n4), .B0(y[19]), .B1(n123), .Y(n121)
         );
  AOI22X1 U98 ( .A0(N89), .A1(n12), .B0(N57), .B1(n5), .Y(n122) );
  CLKINVX1 U99 ( .A(y[19]), .Y(n41) );
  OAI211X1 U100 ( .A0(n81), .A1(n64), .B0(n118), .C0(n119), .Y(N188) );
  AOI32X1 U101 ( .A0(n64), .A1(n39), .A2(n85), .B0(y[20]), .B1(n120), .Y(n118)
         );
  AOI22X1 U102 ( .A0(N90), .A1(n11), .B0(N58), .B1(n5), .Y(n119) );
  CLKINVX1 U103 ( .A(y[20]), .Y(n39) );
  OAI211X1 U104 ( .A0(n14), .A1(n63), .B0(n115), .C0(n116), .Y(N189) );
  AOI32X1 U105 ( .A0(n63), .A1(n38), .A2(n4), .B0(y[21]), .B1(n117), .Y(n115)
         );
  AOI22X1 U106 ( .A0(N91), .A1(n11), .B0(N59), .B1(n5), .Y(n116) );
  CLKINVX1 U107 ( .A(y[21]), .Y(n38) );
  OAI211X1 U108 ( .A0(n81), .A1(n62), .B0(n112), .C0(n113), .Y(N190) );
  AOI32X1 U109 ( .A0(n62), .A1(n37), .A2(n85), .B0(y[22]), .B1(n114), .Y(n112)
         );
  AOI22X1 U110 ( .A0(N92), .A1(n11), .B0(N60), .B1(n5), .Y(n113) );
  CLKINVX1 U111 ( .A(y[22]), .Y(n37) );
  OAI211X1 U112 ( .A0(n14), .A1(n61), .B0(n109), .C0(n110), .Y(N191) );
  AOI32X1 U113 ( .A0(n61), .A1(n36), .A2(n4), .B0(y[23]), .B1(n111), .Y(n109)
         );
  AOI22X1 U114 ( .A0(N93), .A1(n11), .B0(N61), .B1(n5), .Y(n110) );
  CLKINVX1 U115 ( .A(y[23]), .Y(n36) );
  OAI211X1 U116 ( .A0(n81), .A1(n60), .B0(n106), .C0(n107), .Y(N192) );
  AOI32X1 U117 ( .A0(n60), .A1(n35), .A2(n85), .B0(y[24]), .B1(n108), .Y(n106)
         );
  AOI22X1 U118 ( .A0(N94), .A1(n11), .B0(N62), .B1(n5), .Y(n107) );
  CLKINVX1 U119 ( .A(y[24]), .Y(n35) );
  OAI211X1 U120 ( .A0(n14), .A1(n59), .B0(n103), .C0(n104), .Y(N193) );
  AOI32X1 U121 ( .A0(n59), .A1(n34), .A2(n4), .B0(y[25]), .B1(n105), .Y(n103)
         );
  AOI22X1 U122 ( .A0(N95), .A1(n11), .B0(N63), .B1(n5), .Y(n104) );
  CLKINVX1 U123 ( .A(y[25]), .Y(n34) );
  OAI211X1 U124 ( .A0(n81), .A1(n58), .B0(n100), .C0(n101), .Y(N194) );
  AOI32X1 U125 ( .A0(n58), .A1(n33), .A2(n85), .B0(y[26]), .B1(n102), .Y(n100)
         );
  AOI22X1 U126 ( .A0(N96), .A1(n11), .B0(N64), .B1(n5), .Y(n101) );
  CLKINVX1 U127 ( .A(y[26]), .Y(n33) );
  OAI211X1 U128 ( .A0(n14), .A1(n57), .B0(n97), .C0(n98), .Y(N195) );
  AOI32X1 U129 ( .A0(n57), .A1(n32), .A2(n4), .B0(y[27]), .B1(n99), .Y(n97) );
  AOI22X1 U130 ( .A0(N97), .A1(n11), .B0(N65), .B1(n5), .Y(n98) );
  CLKINVX1 U131 ( .A(y[27]), .Y(n32) );
  OAI211X1 U132 ( .A0(n81), .A1(n56), .B0(n94), .C0(n95), .Y(N196) );
  AOI32X1 U133 ( .A0(n56), .A1(n31), .A2(n85), .B0(y[28]), .B1(n96), .Y(n94)
         );
  AOI22X1 U134 ( .A0(N98), .A1(n11), .B0(N66), .B1(n5), .Y(n95) );
  CLKINVX1 U135 ( .A(y[28]), .Y(n31) );
  OAI211X1 U136 ( .A0(n14), .A1(n55), .B0(n91), .C0(n92), .Y(N197) );
  AOI32X1 U137 ( .A0(n55), .A1(n30), .A2(n4), .B0(y[29]), .B1(n93), .Y(n91) );
  AOI22X1 U138 ( .A0(N99), .A1(n11), .B0(N67), .B1(n5), .Y(n92) );
  CLKINVX1 U139 ( .A(y[29]), .Y(n30) );
  OAI211X1 U140 ( .A0(n81), .A1(n54), .B0(n88), .C0(n89), .Y(N198) );
  AOI32X1 U141 ( .A0(n54), .A1(n28), .A2(n85), .B0(y[30]), .B1(n90), .Y(n88)
         );
  AOI22X1 U142 ( .A0(N100), .A1(n11), .B0(N68), .B1(n5), .Y(n89) );
  CLKINVX1 U143 ( .A(y[30]), .Y(n28) );
  NAND4BX2 U144 ( .AN(n4), .B(n184), .C(n8), .D(n181), .Y(N167) );
  NAND3X1 U145 ( .A(ctrl[2]), .B(n52), .C(ctrl[1]), .Y(n184) );
  NOR4X1 U146 ( .A(n52), .B(n19), .C(ctrl[0]), .D(ctrl[1]), .Y(n4) );
  NOR4X1 U147 ( .A(n52), .B(n19), .C(ctrl[0]), .D(ctrl[1]), .Y(n85) );
  CLKINVX1 U148 ( .A(ctrl[2]), .Y(n19) );
  NAND2X1 U149 ( .A(n183), .B(n18), .Y(n87) );
  CLKINVX1 U150 ( .A(ctrl[0]), .Y(n17) );
  CLKINVX1 U151 ( .A(ctrl[1]), .Y(n18) );
  NAND3X1 U152 ( .A(n183), .B(n17), .C(ctrl[1]), .Y(n181) );
  CLKINVX1 U153 ( .A(x[1]), .Y(n187) );
  CLKINVX1 U154 ( .A(x[4]), .Y(n80) );
  CLKINVX1 U155 ( .A(x[5]), .Y(n79) );
  CLKINVX1 U156 ( .A(x[6]), .Y(n78) );
  CLKINVX1 U157 ( .A(x[7]), .Y(n77) );
  CLKINVX1 U158 ( .A(x[14]), .Y(n70) );
  CLKINVX1 U159 ( .A(x[16]), .Y(n68) );
  CLKINVX1 U160 ( .A(x[17]), .Y(n67) );
  CLKINVX1 U161 ( .A(x[22]), .Y(n62) );
  CLKINVX1 U162 ( .A(x[24]), .Y(n60) );
  CLKINVX1 U163 ( .A(x[25]), .Y(n59) );
  CLKINVX1 U164 ( .A(x[30]), .Y(n54) );
  CLKINVX1 U165 ( .A(x[0]), .Y(n188) );
  CLKINVX1 U166 ( .A(x[18]), .Y(n66) );
  CLKINVX1 U167 ( .A(x[26]), .Y(n58) );
  CLKINVX1 U168 ( .A(x[19]), .Y(n65) );
  CLKINVX1 U169 ( .A(x[27]), .Y(n57) );
  CLKINVX1 U170 ( .A(x[21]), .Y(n63) );
  CLKINVX1 U171 ( .A(x[29]), .Y(n55) );
  CLKINVX1 U172 ( .A(x[20]), .Y(n64) );
  CLKINVX1 U173 ( .A(x[28]), .Y(n56) );
  CLKINVX1 U174 ( .A(x[31]), .Y(n53) );
  CLKINVX1 U175 ( .A(x[23]), .Y(n61) );
  CLKBUFX3 U176 ( .A(n84), .Y(n12) );
  CLKBUFX3 U177 ( .A(n84), .Y(n11) );
  CLKBUFX3 U178 ( .A(n81), .Y(n14) );
  NAND3X1 U179 ( .A(n183), .B(n18), .C(ctrl[0]), .Y(n81) );
  CLKBUFX3 U180 ( .A(n84), .Y(n13) );
  OAI211X1 U181 ( .A0(n178), .A1(n51), .B0(n179), .C0(n180), .Y(N168) );
  AOI222XL U182 ( .A0(N38), .A1(n7), .B0(x[0]), .B1(n15), .C0(N70), .C1(n13), 
        .Y(n180) );
  OAI211X1 U183 ( .A0(n14), .A1(n187), .B0(n175), .C0(n176), .Y(N169) );
  AOI22X1 U184 ( .A0(N71), .A1(n13), .B0(N39), .B1(n7), .Y(n176) );
  CLKINVX1 U185 ( .A(y[1]), .Y(n40) );
  OAI211X1 U186 ( .A0(n81), .A1(n76), .B0(n154), .C0(n155), .Y(N176) );
  AOI22X1 U187 ( .A0(N78), .A1(n12), .B0(N46), .B1(n6), .Y(n155) );
  OAI211X1 U188 ( .A0(n14), .A1(n75), .B0(n151), .C0(n152), .Y(N177) );
  AOI22X1 U189 ( .A0(N79), .A1(n12), .B0(N47), .B1(n6), .Y(n152) );
  OAI211X1 U190 ( .A0(n81), .A1(n74), .B0(n148), .C0(n149), .Y(N178) );
  AOI22X1 U191 ( .A0(N80), .A1(n12), .B0(N48), .B1(n6), .Y(n149) );
  OAI211X1 U192 ( .A0(n14), .A1(n73), .B0(n145), .C0(n146), .Y(N179) );
  AOI22X1 U193 ( .A0(N81), .A1(n12), .B0(N49), .B1(n6), .Y(n146) );
  OAI211X1 U194 ( .A0(n81), .A1(n72), .B0(n142), .C0(n143), .Y(N180) );
  AOI22X1 U195 ( .A0(N82), .A1(n12), .B0(N50), .B1(n6), .Y(n143) );
  OAI211X1 U196 ( .A0(n14), .A1(n71), .B0(n139), .C0(n140), .Y(N181) );
  AOI22X1 U197 ( .A0(N83), .A1(n12), .B0(N51), .B1(n6), .Y(n140) );
  OAI211X1 U198 ( .A0(n81), .A1(n70), .B0(n136), .C0(n137), .Y(N182) );
  AOI22X1 U199 ( .A0(N84), .A1(n12), .B0(N52), .B1(n6), .Y(n137) );
  OAI211X1 U200 ( .A0(n14), .A1(n186), .B0(n172), .C0(n173), .Y(N170) );
  AOI32X1 U201 ( .A0(n186), .A1(n29), .A2(n85), .B0(y[2]), .B1(n174), .Y(n172)
         );
  AOI22X1 U202 ( .A0(N72), .A1(n13), .B0(N40), .B1(n7), .Y(n173) );
  CLKINVX1 U203 ( .A(y[2]), .Y(n29) );
  OAI211X1 U204 ( .A0(n81), .A1(n185), .B0(n169), .C0(n170), .Y(N171) );
  AOI32X1 U205 ( .A0(n185), .A1(n26), .A2(n4), .B0(y[3]), .B1(n171), .Y(n169)
         );
  AOI22X1 U206 ( .A0(N73), .A1(n13), .B0(N41), .B1(n7), .Y(n170) );
  CLKINVX1 U207 ( .A(y[3]), .Y(n26) );
  OAI211X1 U208 ( .A0(n14), .A1(n80), .B0(n166), .C0(n167), .Y(N172) );
  AOI32X1 U209 ( .A0(n80), .A1(n25), .A2(n85), .B0(y[4]), .B1(n168), .Y(n166)
         );
  AOI22X1 U210 ( .A0(N74), .A1(n13), .B0(N42), .B1(n7), .Y(n167) );
  CLKINVX1 U211 ( .A(y[4]), .Y(n25) );
  OAI211X1 U212 ( .A0(n81), .A1(n79), .B0(n163), .C0(n164), .Y(N173) );
  AOI32X1 U213 ( .A0(n79), .A1(n24), .A2(n4), .B0(y[5]), .B1(n165), .Y(n163)
         );
  AOI22X1 U214 ( .A0(N75), .A1(n13), .B0(N43), .B1(n7), .Y(n164) );
  CLKINVX1 U215 ( .A(y[5]), .Y(n24) );
  OAI211X1 U216 ( .A0(n14), .A1(n78), .B0(n160), .C0(n161), .Y(N174) );
  AOI22X1 U217 ( .A0(N76), .A1(n13), .B0(N44), .B1(n6), .Y(n161) );
  OAI211X1 U218 ( .A0(n81), .A1(n77), .B0(n157), .C0(n158), .Y(N175) );
  AOI22X1 U219 ( .A0(N77), .A1(n13), .B0(N45), .B1(n6), .Y(n158) );
  NOR2X1 U220 ( .A(ctrl[3]), .B(ctrl[2]), .Y(n183) );
  NOR3X1 U221 ( .A(n17), .B(ctrl[3]), .C(n19), .Y(n182) );
  CLKINVX1 U222 ( .A(ctrl[3]), .Y(n52) );
endmodule


module aluCtrl ( inst, ALUOp, ctrl );
  input [5:0] inst;
  input [1:0] ALUOp;
  output [3:0] ctrl;

  assign ctrl[3] = 1'b0;

  OA21XL U2 ( .A0(inst[0]), .A1(inst[3]), .B0(ALUOp[1]), .Y(ctrl[0]) );
  NAND2X1 U3 ( .A(inst[2]), .B(ALUOp[1]), .Y(ctrl[1]) );
  AO21X1 U4 ( .A0(inst[1]), .A1(ALUOp[1]), .B0(ALUOp[0]), .Y(ctrl[2]) );
endmodule


module control ( inst, inst5_0, RegDst, Jr, Jump, Branch, MemRead, MemToReg, 
        ALUOp, MemWrite, ALUSrc, RegWrite );
  input [5:0] inst;
  input [5:0] inst5_0;
  output [1:0] RegDst;
  output [1:0] MemToReg;
  output [1:0] ALUOp;
  output Jr, Jump, Branch, MemRead, MemWrite, ALUSrc, RegWrite;
  wire   N10, N12, N13, N14, N15, N16, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n1, n2, n3, n4, n5;

  TLATX1 \prev_ALUOp_reg[0]  ( .G(N10), .D(n14), .Q(ALUOp[0]) );
  TLATX1 prev_RegWrite_reg ( .G(N15), .D(N13), .Q(RegWrite) );
  TLATX1 prev_Branch_reg ( .G(N10), .D(n14), .Q(Branch) );
  TLATX1 \prev_RegDst_reg[1]  ( .G(N13), .D(n2), .Q(RegDst[1]) );
  TLATX1 prev_MemWrite_reg ( .G(N15), .D(n13), .Q(MemWrite) );
  TLATX1 \prev_MemToReg_reg[1]  ( .G(N13), .D(n2), .Q(MemToReg[1]) );
  TLATX1 prev_ALUSrc_reg ( .G(N10), .D(n3), .Q(ALUSrc) );
  TLATX1 prev_Jr_reg ( .G(N15), .D(N16), .Q(Jr) );
  TLATX1 \prev_RegDst_reg[0]  ( .G(N13), .D(n15), .Q(RegDst[0]) );
  TLATX1 \prev_ALUOp_reg[1]  ( .G(N10), .D(n15), .Q(ALUOp[1]) );
  TLATX1 prev_MemRead_reg ( .G(N15), .D(n12), .Q(MemRead) );
  TLATX1 prev_Jump_reg ( .G(N15), .D(N14), .Q(Jump) );
  TLATX1 \prev_MemToReg_reg[0]  ( .G(N13), .D(n12), .Q(MemToReg[0]) );
  OR2X1 U3 ( .A(N14), .B(N10), .Y(N15) );
  CLKINVX1 U4 ( .A(n6), .Y(n2) );
  OAI21XL U5 ( .A0(n4), .A1(n8), .B0(n6), .Y(N14) );
  NAND3BX1 U6 ( .AN(n12), .B(n1), .C(n6), .Y(N13) );
  NAND2X1 U7 ( .A(n9), .B(n10), .Y(n6) );
  OR3X2 U8 ( .A(n14), .B(N12), .C(n15), .Y(N10) );
  OR2X1 U9 ( .A(n13), .B(n12), .Y(N12) );
  CLKINVX1 U10 ( .A(n15), .Y(n1) );
  CLKINVX1 U11 ( .A(n11), .Y(n3) );
  NAND3BX1 U12 ( .AN(inst[4]), .B(n10), .C(inst[5]), .Y(n11) );
  NAND3BX1 U13 ( .AN(inst[2]), .B(n9), .C(n5), .Y(n8) );
  NOR3X1 U14 ( .A(inst[4]), .B(inst[5]), .C(inst[3]), .Y(n9) );
  NOR4BX1 U15 ( .AN(inst5_0[3]), .B(n7), .C(inst5_0[0]), .D(n1), .Y(N16) );
  OR4X1 U16 ( .A(inst5_0[2]), .B(inst5_0[1]), .C(inst5_0[5]), .D(inst5_0[4]), 
        .Y(n7) );
  NOR3X1 U17 ( .A(n5), .B(inst[2]), .C(n4), .Y(n10) );
  NOR2X1 U18 ( .A(n8), .B(inst[1]), .Y(n15) );
  NOR2BX1 U19 ( .AN(inst[3]), .B(n11), .Y(n13) );
  NOR2X1 U20 ( .A(n11), .B(inst[3]), .Y(n12) );
  AND4X1 U21 ( .A(inst[2]), .B(n9), .C(n5), .D(n4), .Y(n14) );
  CLKINVX1 U22 ( .A(inst[1]), .Y(n4) );
  CLKINVX1 U23 ( .A(inst[0]), .Y(n5) );
endmodule


module SingleCycle_MIPS_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30;

  XOR2X1 U1 ( .A(A[29]), .B(n24), .Y(SUM[29]) );
  XOR2X1 U2 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  XOR2X1 U3 ( .A(A[5]), .B(n2), .Y(SUM[5]) );
  XOR2X1 U4 ( .A(A[6]), .B(n3), .Y(SUM[6]) );
  XOR2X1 U5 ( .A(A[7]), .B(n4), .Y(SUM[7]) );
  XOR2X1 U6 ( .A(A[8]), .B(n5), .Y(SUM[8]) );
  XOR2X1 U7 ( .A(A[9]), .B(n6), .Y(SUM[9]) );
  XOR2X1 U8 ( .A(A[10]), .B(n7), .Y(SUM[10]) );
  XOR2X1 U9 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  XOR2X1 U10 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2X1 U11 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  CLKINVX1 U12 ( .A(A[2]), .Y(SUM[2]) );
  AND2X2 U13 ( .A(A[3]), .B(A[2]), .Y(n1) );
  AND2X2 U14 ( .A(A[4]), .B(n1), .Y(n2) );
  AND2X2 U15 ( .A(A[5]), .B(n2), .Y(n3) );
  AND2X2 U16 ( .A(A[6]), .B(n3), .Y(n4) );
  AND2X2 U17 ( .A(A[7]), .B(n4), .Y(n5) );
  AND2X2 U18 ( .A(A[8]), .B(n5), .Y(n6) );
  AND2X2 U19 ( .A(A[9]), .B(n6), .Y(n7) );
  AND2X2 U20 ( .A(A[10]), .B(n7), .Y(n8) );
  AND2X2 U21 ( .A(A[11]), .B(n8), .Y(n9) );
  XNOR2X1 U22 ( .A(A[31]), .B(n30), .Y(SUM[31]) );
  NAND2X1 U23 ( .A(A[30]), .B(n25), .Y(n30) );
  XOR2X1 U24 ( .A(A[28]), .B(n23), .Y(SUM[28]) );
  XOR2X1 U25 ( .A(A[13]), .B(n26), .Y(SUM[13]) );
  XOR2X1 U26 ( .A(A[14]), .B(n27), .Y(SUM[14]) );
  XOR2X1 U27 ( .A(A[15]), .B(n10), .Y(SUM[15]) );
  XOR2X1 U28 ( .A(A[16]), .B(n11), .Y(SUM[16]) );
  XOR2X1 U29 ( .A(A[17]), .B(n12), .Y(SUM[17]) );
  XOR2X1 U30 ( .A(A[18]), .B(n13), .Y(SUM[18]) );
  XOR2X1 U31 ( .A(A[19]), .B(n14), .Y(SUM[19]) );
  XOR2X1 U32 ( .A(A[20]), .B(n15), .Y(SUM[20]) );
  XOR2X1 U33 ( .A(A[21]), .B(n16), .Y(SUM[21]) );
  XOR2X1 U34 ( .A(A[22]), .B(n17), .Y(SUM[22]) );
  XOR2X1 U35 ( .A(A[23]), .B(n18), .Y(SUM[23]) );
  XOR2X1 U36 ( .A(A[24]), .B(n19), .Y(SUM[24]) );
  XOR2X1 U37 ( .A(A[25]), .B(n20), .Y(SUM[25]) );
  XOR2X1 U38 ( .A(A[26]), .B(n21), .Y(SUM[26]) );
  XOR2X1 U39 ( .A(A[27]), .B(n22), .Y(SUM[27]) );
  AND2X2 U40 ( .A(A[14]), .B(n27), .Y(n10) );
  AND2X2 U41 ( .A(A[15]), .B(n10), .Y(n11) );
  AND2X2 U42 ( .A(A[16]), .B(n11), .Y(n12) );
  AND2X2 U43 ( .A(A[17]), .B(n12), .Y(n13) );
  AND2X2 U44 ( .A(A[18]), .B(n13), .Y(n14) );
  AND2X2 U45 ( .A(A[19]), .B(n14), .Y(n15) );
  AND2X2 U46 ( .A(A[20]), .B(n15), .Y(n16) );
  AND2X2 U47 ( .A(A[21]), .B(n16), .Y(n17) );
  AND2X2 U48 ( .A(A[22]), .B(n17), .Y(n18) );
  AND2X2 U49 ( .A(A[23]), .B(n18), .Y(n19) );
  AND2X2 U50 ( .A(A[24]), .B(n19), .Y(n20) );
  AND2X2 U51 ( .A(A[25]), .B(n20), .Y(n21) );
  AND2X2 U52 ( .A(A[26]), .B(n21), .Y(n22) );
  AND2X2 U53 ( .A(A[27]), .B(n22), .Y(n23) );
  AND2X2 U54 ( .A(A[28]), .B(n23), .Y(n24) );
  AND2X2 U55 ( .A(A[29]), .B(n24), .Y(n25) );
  AND2X2 U56 ( .A(A[12]), .B(n9), .Y(n26) );
  AND2X2 U57 ( .A(A[13]), .B(n26), .Y(n27) );
  XOR2X1 U58 ( .A(A[30]), .B(n25), .Y(SUM[30]) );
  CLKBUFX3 U59 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U60 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SingleCycle_MIPS_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2XL U2 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U3 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U4 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SingleCycle_MIPS ( clk, rst_n, IR_addr, IR, RF_writedata, ReadDataMem, 
        CEN, WEN, A, ReadData2, OEN );
  output [31:0] IR_addr;
  input [31:0] IR;
  output [31:0] RF_writedata;
  input [31:0] ReadDataMem;
  output [6:0] A;
  output [31:0] ReadData2;
  input clk, rst_n;
  output CEN, WEN, OEN;
  wire   RegWrite, zero, ALUResult_1, ALUResult_0, Jump, Jr, Branch, MemRead,
         MemWrite, ALUSrc, n67, n68, n69, n70, n71, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n85, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, N57, N42, N41, N40, N39, N38, N37, N36,
         N35, N34, N33, N32, N31, N30, N29, N28, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209;
  wire   [31:0] ReadData1;
  wire   [3:0] ctrl;
  wire   [31:0] y;
  wire   [31:9] ALUResult;
  wire   [1:0] ALUOp;
  wire   [1:0] RegDst;
  wire   [1:0] MemToReg;
  wire   [31:0] next_address;
  wire   [31:0] muxres1;
  wire   [31:0] muxres3;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign OEN = 1'b0;

  register register ( .clk(clk), .rst_n(n179), .RegWrite(RegWrite), .ReadReg1(
        {IR[25], n178, IR[23], n177, n176}), .ReadReg2({IR[20], n175, n174, 
        n173, n172}), .WriteReg({n67, n68, n69, n70, n71}), .WriteData(
        RF_writedata), .ReadData1(ReadData1), .ReadData2(ReadData2) );
  alu alu ( .ctrl({1'b0, ctrl[2:0]}), .x(ReadData1), .y(y), .zero(zero), .out(
        {ALUResult, A, ALUResult_1, ALUResult_0}) );
  aluCtrl aluCtrl ( .inst(IR[5:0]), .ALUOp(ALUOp), .ctrl({
        SYNOPSYS_UNCONNECTED__0, ctrl[2:0]}) );
  control control ( .inst(IR[31:26]), .inst5_0(IR[5:0]), .RegDst(RegDst), .Jr(
        Jr), .Jump(Jump), .Branch(Branch), .MemRead(MemRead), .MemToReg(
        MemToReg), .ALUOp(ALUOp), .MemWrite(MemWrite), .ALUSrc(ALUSrc), 
        .RegWrite(RegWrite) );
  SingleCycle_MIPS_DW01_add_0 add_106 ( .A(IR_addr), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(next_address) );
  SingleCycle_MIPS_DW01_add_1 add_110_aco ( .A(next_address), .B({n165, n164, 
        n165, n164, n165, n164, n165, n164, n165, n164, n165, n164, n165, n164, 
        n164, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, 1'b0, 1'b0}), .CI(1'b0), .SUM(muxres1) );
  DFFRX1 \reg_IR_addr_reg[0]  ( .D(muxres3[0]), .CK(clk), .RN(n179), .Q(
        IR_addr[0]) );
  DFFRX1 \reg_IR_addr_reg[1]  ( .D(muxres3[1]), .CK(clk), .RN(n179), .Q(
        IR_addr[1]) );
  DFFRX1 \reg_IR_addr_reg[31]  ( .D(n181), .CK(clk), .RN(n179), .Q(IR_addr[31]) );
  DFFRX1 \reg_IR_addr_reg[23]  ( .D(n186), .CK(clk), .RN(n179), .Q(IR_addr[23]) );
  DFFRX1 \reg_IR_addr_reg[24]  ( .D(n185), .CK(clk), .RN(n179), .Q(IR_addr[24]) );
  DFFRX1 \reg_IR_addr_reg[25]  ( .D(n184), .CK(clk), .RN(n179), .Q(IR_addr[25]) );
  DFFRX1 \reg_IR_addr_reg[26]  ( .D(n183), .CK(clk), .RN(n179), .Q(IR_addr[26]) );
  DFFRX1 \reg_IR_addr_reg[27]  ( .D(n182), .CK(clk), .RN(n179), .Q(IR_addr[27]) );
  DFFRX1 \reg_IR_addr_reg[28]  ( .D(n146), .CK(clk), .RN(n179), .Q(IR_addr[28]) );
  DFFRX1 \reg_IR_addr_reg[29]  ( .D(n147), .CK(clk), .RN(n179), .Q(IR_addr[29]) );
  DFFRX1 \reg_IR_addr_reg[14]  ( .D(n195), .CK(clk), .RN(n179), .Q(IR_addr[14]) );
  DFFRX1 \reg_IR_addr_reg[15]  ( .D(n194), .CK(clk), .RN(n179), .Q(IR_addr[15]) );
  DFFRX1 \reg_IR_addr_reg[16]  ( .D(n193), .CK(clk), .RN(n179), .Q(IR_addr[16]) );
  DFFRX1 \reg_IR_addr_reg[17]  ( .D(n192), .CK(clk), .RN(n179), .Q(IR_addr[17]) );
  DFFRX1 \reg_IR_addr_reg[18]  ( .D(n191), .CK(clk), .RN(n179), .Q(IR_addr[18]) );
  DFFRX1 \reg_IR_addr_reg[19]  ( .D(n190), .CK(clk), .RN(n179), .Q(IR_addr[19]) );
  DFFRX1 \reg_IR_addr_reg[20]  ( .D(n189), .CK(clk), .RN(n179), .Q(IR_addr[20]) );
  DFFRX1 \reg_IR_addr_reg[21]  ( .D(n188), .CK(clk), .RN(n179), .Q(IR_addr[21]) );
  DFFRX1 \reg_IR_addr_reg[22]  ( .D(n187), .CK(clk), .RN(n179), .Q(IR_addr[22]) );
  DFFRX1 \reg_IR_addr_reg[5]  ( .D(n204), .CK(clk), .RN(n179), .Q(IR_addr[5])
         );
  DFFRX1 \reg_IR_addr_reg[6]  ( .D(n203), .CK(clk), .RN(n179), .Q(IR_addr[6])
         );
  DFFRX1 \reg_IR_addr_reg[7]  ( .D(n202), .CK(clk), .RN(n179), .Q(IR_addr[7])
         );
  DFFRX1 \reg_IR_addr_reg[8]  ( .D(n201), .CK(clk), .RN(n179), .Q(IR_addr[8])
         );
  DFFRX1 \reg_IR_addr_reg[9]  ( .D(n200), .CK(clk), .RN(n179), .Q(IR_addr[9])
         );
  DFFRX1 \reg_IR_addr_reg[10]  ( .D(n199), .CK(clk), .RN(n179), .Q(IR_addr[10]) );
  DFFRX1 \reg_IR_addr_reg[11]  ( .D(n198), .CK(clk), .RN(n179), .Q(IR_addr[11]) );
  DFFRX1 \reg_IR_addr_reg[12]  ( .D(n197), .CK(clk), .RN(n179), .Q(IR_addr[12]) );
  DFFRX1 \reg_IR_addr_reg[13]  ( .D(n196), .CK(clk), .RN(n179), .Q(IR_addr[13]) );
  DFFRX1 \reg_IR_addr_reg[3]  ( .D(n206), .CK(clk), .RN(n179), .Q(IR_addr[3])
         );
  DFFRX1 \reg_IR_addr_reg[4]  ( .D(n205), .CK(clk), .RN(n179), .Q(IR_addr[4])
         );
  DFFRX1 \reg_IR_addr_reg[2]  ( .D(n207), .CK(clk), .RN(n179), .Q(IR_addr[2])
         );
  TLATNX1 prev_WEN_reg ( .D(MemRead), .GN(CEN), .Q(WEN) );
  DFFRX1 \reg_IR_addr_reg[30]  ( .D(n154), .CK(clk), .RN(n179), .Q(IR_addr[30]) );
  NOR2X1 U214 ( .A(MemToReg[0]), .B(n170), .Y(n112) );
  NOR2X1 U215 ( .A(n171), .B(Jump), .Y(n76) );
  AOI222X1 U216 ( .A0(ReadData1[31]), .A1(n171), .B0(next_address[31]), .B1(
        n169), .C0(muxres1[31]), .C1(n76), .Y(n83) );
  OR3X2 U217 ( .A(n148), .B(n149), .C(n150), .Y(n146) );
  NAND3X1 U218 ( .A(n151), .B(n152), .C(n153), .Y(n147) );
  NAND2X1 U219 ( .A(n158), .B(n159), .Y(y[0]) );
  NAND2X1 U220 ( .A(ReadData2[0]), .B(n209), .Y(n159) );
  AND2X2 U221 ( .A(next_address[28]), .B(n169), .Y(n149) );
  AND2X2 U222 ( .A(muxres1[28]), .B(n76), .Y(n150) );
  INVXL U223 ( .A(n88), .Y(n182) );
  AND2X2 U224 ( .A(ReadData1[28]), .B(n171), .Y(n148) );
  INVXL U225 ( .A(n83), .Y(n181) );
  NAND2XL U226 ( .A(muxres1[29]), .B(n76), .Y(n153) );
  NAND2XL U227 ( .A(zero), .B(Branch), .Y(n160) );
  NAND2X1 U228 ( .A(muxres1[30]), .B(n76), .Y(n157) );
  AOI222XL U229 ( .A0(ReadData1[26]), .A1(n171), .B0(n178), .B1(n75), .C0(
        muxres1[26]), .C1(n76), .Y(n89) );
  AO22X1 U230 ( .A0(n163), .A1(IR[4]), .B0(ReadData2[4]), .B1(n209), .Y(y[4])
         );
  AO22X1 U231 ( .A0(n163), .A1(IR[5]), .B0(ReadData2[5]), .B1(n209), .Y(y[5])
         );
  AO22X1 U232 ( .A0(n163), .A1(IR[1]), .B0(ReadData2[1]), .B1(n209), .Y(y[1])
         );
  AO22X1 U233 ( .A0(n163), .A1(IR[2]), .B0(ReadData2[2]), .B1(n209), .Y(y[2])
         );
  AO22X1 U234 ( .A0(n163), .A1(IR[3]), .B0(ReadData2[3]), .B1(n209), .Y(y[3])
         );
  NAND2X1 U235 ( .A(zero), .B(Branch), .Y(n162) );
  NAND2X1 U236 ( .A(ReadData1[29]), .B(n171), .Y(n151) );
  NAND2X1 U237 ( .A(next_address[29]), .B(n75), .Y(n152) );
  NAND3X1 U238 ( .A(n155), .B(n156), .C(n157), .Y(n154) );
  AOI222XL U239 ( .A0(next_address[0]), .A1(n170), .B0(ALUResult_0), .B1(n112), 
        .C0(ReadDataMem[0]), .C1(n166), .Y(n144) );
  AOI222XL U240 ( .A0(next_address[1]), .A1(n170), .B0(ALUResult_1), .B1(n112), 
        .C0(ReadDataMem[1]), .C1(n113), .Y(n133) );
  AOI222XL U241 ( .A0(next_address[2]), .A1(n170), .B0(A[0]), .B1(n112), .C0(
        ReadDataMem[2]), .C1(n167), .Y(n122) );
  AOI222XL U242 ( .A0(next_address[3]), .A1(n170), .B0(A[1]), .B1(n112), .C0(
        ReadDataMem[3]), .C1(n167), .Y(n119) );
  AOI222XL U243 ( .A0(next_address[4]), .A1(n170), .B0(A[2]), .B1(n112), .C0(
        ReadDataMem[4]), .C1(n113), .Y(n118) );
  AOI222XL U244 ( .A0(next_address[5]), .A1(n170), .B0(A[3]), .B1(n112), .C0(
        ReadDataMem[5]), .C1(n166), .Y(n117) );
  AOI222XL U245 ( .A0(next_address[6]), .A1(n170), .B0(A[4]), .B1(n112), .C0(
        ReadDataMem[6]), .C1(n167), .Y(n116) );
  AOI222XL U246 ( .A0(next_address[7]), .A1(n170), .B0(A[5]), .B1(n112), .C0(
        ReadDataMem[7]), .C1(n113), .Y(n115) );
  AOI222XL U247 ( .A0(next_address[8]), .A1(n170), .B0(A[6]), .B1(n112), .C0(
        ReadDataMem[8]), .C1(n166), .Y(n114) );
  AOI222XL U248 ( .A0(next_address[9]), .A1(n170), .B0(ALUResult[9]), .B1(n112), .C0(ReadDataMem[9]), .C1(n167), .Y(n111) );
  AOI222XL U249 ( .A0(next_address[10]), .A1(n170), .B0(ALUResult[10]), .B1(
        n112), .C0(ReadDataMem[10]), .C1(n167), .Y(n143) );
  AOI222XL U250 ( .A0(next_address[11]), .A1(n170), .B0(ALUResult[11]), .B1(
        n112), .C0(ReadDataMem[11]), .C1(n113), .Y(n142) );
  AOI222XL U251 ( .A0(next_address[12]), .A1(n170), .B0(ALUResult[12]), .B1(
        n112), .C0(ReadDataMem[12]), .C1(n166), .Y(n141) );
  AOI222XL U252 ( .A0(next_address[13]), .A1(n170), .B0(ALUResult[13]), .B1(
        n112), .C0(ReadDataMem[13]), .C1(n167), .Y(n140) );
  AOI222XL U253 ( .A0(next_address[14]), .A1(n170), .B0(ALUResult[14]), .B1(
        n112), .C0(ReadDataMem[14]), .C1(n113), .Y(n139) );
  AOI222XL U254 ( .A0(next_address[15]), .A1(n170), .B0(ALUResult[15]), .B1(
        n112), .C0(ReadDataMem[15]), .C1(n166), .Y(n138) );
  AOI222XL U255 ( .A0(next_address[16]), .A1(n170), .B0(ALUResult[16]), .B1(
        n112), .C0(ReadDataMem[16]), .C1(n167), .Y(n137) );
  AOI222XL U256 ( .A0(next_address[17]), .A1(n170), .B0(ALUResult[17]), .B1(
        n112), .C0(ReadDataMem[17]), .C1(n113), .Y(n136) );
  AOI222XL U257 ( .A0(next_address[18]), .A1(n170), .B0(ALUResult[18]), .B1(
        n112), .C0(ReadDataMem[18]), .C1(n166), .Y(n135) );
  AOI222XL U258 ( .A0(next_address[19]), .A1(n170), .B0(ALUResult[19]), .B1(
        n112), .C0(ReadDataMem[19]), .C1(n167), .Y(n134) );
  AOI222XL U259 ( .A0(next_address[20]), .A1(n170), .B0(ALUResult[20]), .B1(
        n112), .C0(ReadDataMem[20]), .C1(n166), .Y(n132) );
  AOI222XL U260 ( .A0(next_address[21]), .A1(n170), .B0(ALUResult[21]), .B1(
        n112), .C0(ReadDataMem[21]), .C1(n167), .Y(n131) );
  AOI222XL U261 ( .A0(next_address[22]), .A1(n170), .B0(ALUResult[22]), .B1(
        n112), .C0(ReadDataMem[22]), .C1(n113), .Y(n130) );
  AOI222XL U262 ( .A0(next_address[23]), .A1(n170), .B0(ALUResult[23]), .B1(
        n112), .C0(ReadDataMem[23]), .C1(n166), .Y(n129) );
  AOI222XL U263 ( .A0(next_address[24]), .A1(n170), .B0(ALUResult[24]), .B1(
        n112), .C0(ReadDataMem[24]), .C1(n167), .Y(n128) );
  AOI222XL U264 ( .A0(next_address[25]), .A1(n170), .B0(ALUResult[25]), .B1(
        n112), .C0(ReadDataMem[25]), .C1(n113), .Y(n127) );
  AOI222XL U265 ( .A0(next_address[26]), .A1(n170), .B0(ALUResult[26]), .B1(
        n112), .C0(ReadDataMem[26]), .C1(n166), .Y(n126) );
  AOI222XL U266 ( .A0(next_address[27]), .A1(n170), .B0(ALUResult[27]), .B1(
        n112), .C0(ReadDataMem[27]), .C1(n167), .Y(n125) );
  AOI222XL U267 ( .A0(n170), .A1(next_address[28]), .B0(ALUResult[28]), .B1(
        n112), .C0(ReadDataMem[28]), .C1(n113), .Y(n124) );
  AOI222XL U268 ( .A0(n170), .A1(next_address[29]), .B0(ALUResult[29]), .B1(
        n112), .C0(ReadDataMem[29]), .C1(n166), .Y(n123) );
  AOI222XL U269 ( .A0(n170), .A1(next_address[30]), .B0(ALUResult[30]), .B1(
        n112), .C0(ReadDataMem[30]), .C1(n113), .Y(n121) );
  AOI222XL U270 ( .A0(n170), .A1(next_address[31]), .B0(ALUResult[31]), .B1(
        n112), .C0(ReadDataMem[31]), .C1(n166), .Y(n120) );
  NAND2X1 U271 ( .A(IR[15]), .B(n163), .Y(n73) );
  CLKINVX1 U272 ( .A(n108), .Y(n69) );
  CLKINVX1 U273 ( .A(n110), .Y(n71) );
  CLKINVX1 U274 ( .A(n109), .Y(n70) );
  CLKBUFX3 U275 ( .A(ALUSrc), .Y(n163) );
  NAND2X1 U276 ( .A(ReadData1[30]), .B(n171), .Y(n155) );
  NAND2X1 U277 ( .A(next_address[30]), .B(n168), .Y(n156) );
  NAND2X1 U278 ( .A(n163), .B(IR[0]), .Y(n158) );
  NAND2XL U279 ( .A(zero), .B(Branch), .Y(n161) );
  CLKINVX1 U280 ( .A(n89), .Y(n183) );
  OAI2BB1X1 U281 ( .A0N(ReadData2[18]), .A1N(n209), .B0(n73), .Y(y[18]) );
  OAI2BB1X1 U282 ( .A0N(ReadData2[19]), .A1N(n209), .B0(n73), .Y(y[19]) );
  OAI2BB1X1 U283 ( .A0N(ReadData2[20]), .A1N(n209), .B0(n73), .Y(y[20]) );
  OAI2BB1X1 U284 ( .A0N(ReadData2[21]), .A1N(n209), .B0(n73), .Y(y[21]) );
  OAI2BB1X1 U285 ( .A0N(ReadData2[15]), .A1N(n209), .B0(n73), .Y(y[15]) );
  OAI2BB1X1 U286 ( .A0N(ReadData2[16]), .A1N(n209), .B0(n73), .Y(y[16]) );
  OAI2BB1X1 U287 ( .A0N(ReadData2[17]), .A1N(n209), .B0(n73), .Y(y[17]) );
  OAI2BB1X1 U288 ( .A0N(ReadData2[22]), .A1N(n209), .B0(n73), .Y(y[22]) );
  CLKBUFX3 U289 ( .A(N57), .Y(n164) );
  CLKBUFX3 U290 ( .A(N57), .Y(n165) );
  CLKINVX1 U291 ( .A(n91), .Y(n185) );
  AOI222XL U292 ( .A0(ReadData1[24]), .A1(n171), .B0(n177), .B1(n168), .C0(
        muxres1[24]), .C1(n76), .Y(n91) );
  CLKINVX1 U293 ( .A(n92), .Y(n186) );
  AOI222XL U294 ( .A0(ReadData1[23]), .A1(n171), .B0(n176), .B1(n75), .C0(
        muxres1[23]), .C1(n76), .Y(n92) );
  CLKINVX1 U295 ( .A(n94), .Y(n188) );
  AOI222XL U296 ( .A0(ReadData1[21]), .A1(n171), .B0(n175), .B1(n168), .C0(
        muxres1[21]), .C1(n76), .Y(n94) );
  CLKINVX1 U297 ( .A(n95), .Y(n189) );
  AOI222XL U298 ( .A0(ReadData1[20]), .A1(n171), .B0(n174), .B1(n75), .C0(
        muxres1[20]), .C1(n76), .Y(n95) );
  CLKINVX1 U299 ( .A(n96), .Y(n190) );
  AOI222XL U300 ( .A0(ReadData1[19]), .A1(n171), .B0(n173), .B1(n169), .C0(
        muxres1[19]), .C1(n76), .Y(n96) );
  CLKINVX1 U301 ( .A(n97), .Y(n191) );
  AOI222XL U302 ( .A0(ReadData1[18]), .A1(n171), .B0(n172), .B1(n168), .C0(
        muxres1[18]), .C1(n76), .Y(n97) );
  CLKINVX1 U303 ( .A(n124), .Y(RF_writedata[28]) );
  CLKINVX1 U304 ( .A(n123), .Y(RF_writedata[29]) );
  CLKINVX1 U305 ( .A(n121), .Y(RF_writedata[30]) );
  CLKINVX1 U306 ( .A(n120), .Y(RF_writedata[31]) );
  CLKINVX1 U307 ( .A(n144), .Y(RF_writedata[0]) );
  CLKINVX1 U308 ( .A(n133), .Y(RF_writedata[1]) );
  CLKINVX1 U309 ( .A(n122), .Y(RF_writedata[2]) );
  CLKINVX1 U310 ( .A(n119), .Y(RF_writedata[3]) );
  CLKINVX1 U311 ( .A(n118), .Y(RF_writedata[4]) );
  CLKINVX1 U312 ( .A(n117), .Y(RF_writedata[5]) );
  CLKINVX1 U313 ( .A(n116), .Y(RF_writedata[6]) );
  CLKINVX1 U314 ( .A(n115), .Y(RF_writedata[7]) );
  CLKINVX1 U315 ( .A(n114), .Y(RF_writedata[8]) );
  CLKINVX1 U316 ( .A(n111), .Y(RF_writedata[9]) );
  CLKINVX1 U317 ( .A(n143), .Y(RF_writedata[10]) );
  CLKINVX1 U318 ( .A(n142), .Y(RF_writedata[11]) );
  CLKINVX1 U319 ( .A(n141), .Y(RF_writedata[12]) );
  CLKINVX1 U320 ( .A(n140), .Y(RF_writedata[13]) );
  CLKINVX1 U321 ( .A(n139), .Y(RF_writedata[14]) );
  CLKINVX1 U322 ( .A(n138), .Y(RF_writedata[15]) );
  CLKINVX1 U323 ( .A(n137), .Y(RF_writedata[16]) );
  CLKINVX1 U324 ( .A(n136), .Y(RF_writedata[17]) );
  CLKINVX1 U325 ( .A(n135), .Y(RF_writedata[18]) );
  CLKINVX1 U326 ( .A(n134), .Y(RF_writedata[19]) );
  CLKINVX1 U327 ( .A(n132), .Y(RF_writedata[20]) );
  CLKINVX1 U328 ( .A(n131), .Y(RF_writedata[21]) );
  CLKINVX1 U329 ( .A(n130), .Y(RF_writedata[22]) );
  CLKINVX1 U330 ( .A(n129), .Y(RF_writedata[23]) );
  CLKINVX1 U331 ( .A(n128), .Y(RF_writedata[24]) );
  CLKINVX1 U332 ( .A(n127), .Y(RF_writedata[25]) );
  CLKINVX1 U333 ( .A(n126), .Y(RF_writedata[26]) );
  CLKINVX1 U334 ( .A(n125), .Y(RF_writedata[27]) );
  OAI2BB1X1 U335 ( .A0N(ReadData2[31]), .A1N(n209), .B0(n73), .Y(y[31]) );
  OAI2BB1X1 U336 ( .A0N(ReadData2[26]), .A1N(n209), .B0(n73), .Y(y[26]) );
  OAI2BB1X1 U337 ( .A0N(ReadData2[27]), .A1N(n209), .B0(n73), .Y(y[27]) );
  OAI2BB1X1 U338 ( .A0N(ReadData2[28]), .A1N(n209), .B0(n73), .Y(y[28]) );
  OAI2BB1X1 U339 ( .A0N(ReadData2[29]), .A1N(n209), .B0(n73), .Y(y[29]) );
  OAI2BB1X1 U340 ( .A0N(ReadData2[23]), .A1N(n209), .B0(n73), .Y(y[23]) );
  OAI2BB1X1 U341 ( .A0N(ReadData2[24]), .A1N(n209), .B0(n73), .Y(y[24]) );
  OAI2BB1X1 U342 ( .A0N(ReadData2[25]), .A1N(n209), .B0(n73), .Y(y[25]) );
  OAI2BB1X1 U343 ( .A0N(ReadData2[30]), .A1N(n209), .B0(n73), .Y(y[30]) );
  AO22X1 U344 ( .A0(ReadData1[0]), .A1(n171), .B0(muxres1[0]), .B1(n76), .Y(
        muxres3[0]) );
  AO22X1 U345 ( .A0(ReadData1[1]), .A1(n171), .B0(muxres1[1]), .B1(n76), .Y(
        muxres3[1]) );
  CLKINVX1 U346 ( .A(n163), .Y(n209) );
  AO22X1 U347 ( .A0(n163), .A1(IR[8]), .B0(ReadData2[8]), .B1(n209), .Y(y[8])
         );
  AO22X1 U348 ( .A0(n163), .A1(IR[6]), .B0(ReadData2[6]), .B1(n209), .Y(y[6])
         );
  AO22X1 U349 ( .A0(n163), .A1(IR[7]), .B0(ReadData2[7]), .B1(n209), .Y(y[7])
         );
  AOI222XL U350 ( .A0(ReadData1[27]), .A1(n171), .B0(IR[25]), .B1(n168), .C0(
        muxres1[27]), .C1(n76), .Y(n88) );
  CLKINVX1 U351 ( .A(n90), .Y(n184) );
  AOI222XL U352 ( .A0(ReadData1[25]), .A1(n171), .B0(IR[23]), .B1(n169), .C0(
        muxres1[25]), .C1(n76), .Y(n90) );
  AO22X1 U353 ( .A0(n163), .A1(IR[9]), .B0(ReadData2[9]), .B1(n209), .Y(y[9])
         );
  AO22X1 U354 ( .A0(n163), .A1(IR[10]), .B0(ReadData2[10]), .B1(n209), .Y(
        y[10]) );
  AO22X1 U355 ( .A0(n163), .A1(IR[11]), .B0(ReadData2[11]), .B1(n209), .Y(
        y[11]) );
  AO22X1 U356 ( .A0(n163), .A1(IR[12]), .B0(ReadData2[12]), .B1(n209), .Y(
        y[12]) );
  AO22X1 U357 ( .A0(n163), .A1(IR[13]), .B0(ReadData2[13]), .B1(n209), .Y(
        y[13]) );
  AO22X1 U358 ( .A0(n163), .A1(IR[14]), .B0(ReadData2[14]), .B1(n209), .Y(
        y[14]) );
  NOR2X1 U359 ( .A(n160), .B(n180), .Y(N57) );
  CLKINVX1 U360 ( .A(IR[15]), .Y(n180) );
  CLKINVX1 U361 ( .A(n93), .Y(n187) );
  AOI222XL U362 ( .A0(ReadData1[22]), .A1(n171), .B0(IR[20]), .B1(n169), .C0(
        muxres1[22]), .C1(n76), .Y(n93) );
  CLKINVX1 U363 ( .A(n98), .Y(n192) );
  AOI222XL U364 ( .A0(ReadData1[17]), .A1(n171), .B0(n168), .B1(IR[15]), .C0(
        muxres1[17]), .C1(n76), .Y(n98) );
  CLKINVX1 U365 ( .A(n99), .Y(n193) );
  AOI222XL U366 ( .A0(ReadData1[16]), .A1(n171), .B0(n75), .B1(IR[14]), .C0(
        muxres1[16]), .C1(n76), .Y(n99) );
  CLKINVX1 U367 ( .A(n100), .Y(n194) );
  AOI222XL U368 ( .A0(ReadData1[15]), .A1(n171), .B0(n169), .B1(IR[13]), .C0(
        muxres1[15]), .C1(n76), .Y(n100) );
  CLKINVX1 U369 ( .A(n101), .Y(n195) );
  AOI222XL U370 ( .A0(ReadData1[14]), .A1(n171), .B0(n168), .B1(IR[12]), .C0(
        muxres1[14]), .C1(n76), .Y(n101) );
  CLKINVX1 U371 ( .A(n102), .Y(n196) );
  AOI222XL U372 ( .A0(ReadData1[13]), .A1(n171), .B0(n75), .B1(IR[11]), .C0(
        muxres1[13]), .C1(n76), .Y(n102) );
  CLKINVX1 U373 ( .A(n85), .Y(n207) );
  AOI222XL U374 ( .A0(ReadData1[2]), .A1(n171), .B0(n169), .B1(IR[0]), .C0(
        muxres1[2]), .C1(n76), .Y(n85) );
  CLKINVX1 U375 ( .A(n103), .Y(n197) );
  AOI222XL U376 ( .A0(ReadData1[12]), .A1(n171), .B0(n169), .B1(IR[10]), .C0(
        muxres1[12]), .C1(n76), .Y(n103) );
  CLKINVX1 U377 ( .A(n104), .Y(n198) );
  AOI222XL U378 ( .A0(ReadData1[11]), .A1(n171), .B0(n168), .B1(IR[9]), .C0(
        muxres1[11]), .C1(n76), .Y(n104) );
  CLKINVX1 U379 ( .A(n105), .Y(n199) );
  AOI222XL U380 ( .A0(ReadData1[10]), .A1(n171), .B0(n75), .B1(IR[8]), .C0(
        muxres1[10]), .C1(n76), .Y(n105) );
  CLKINVX1 U381 ( .A(n74), .Y(n200) );
  AOI222XL U382 ( .A0(ReadData1[9]), .A1(n171), .B0(n75), .B1(IR[7]), .C0(
        muxres1[9]), .C1(n76), .Y(n74) );
  CLKINVX1 U383 ( .A(n77), .Y(n201) );
  AOI222XL U384 ( .A0(ReadData1[8]), .A1(n171), .B0(n169), .B1(IR[6]), .C0(
        muxres1[8]), .C1(n76), .Y(n77) );
  CLKINVX1 U385 ( .A(n78), .Y(n202) );
  AOI222XL U386 ( .A0(ReadData1[7]), .A1(n171), .B0(n168), .B1(IR[5]), .C0(
        muxres1[7]), .C1(n76), .Y(n78) );
  CLKINVX1 U387 ( .A(n79), .Y(n203) );
  AOI222XL U388 ( .A0(ReadData1[6]), .A1(n171), .B0(n75), .B1(IR[4]), .C0(
        muxres1[6]), .C1(n76), .Y(n79) );
  CLKINVX1 U389 ( .A(n80), .Y(n204) );
  AOI222XL U390 ( .A0(ReadData1[5]), .A1(n171), .B0(n169), .B1(IR[3]), .C0(
        muxres1[5]), .C1(n76), .Y(n80) );
  CLKINVX1 U391 ( .A(n81), .Y(n205) );
  AOI222XL U392 ( .A0(ReadData1[4]), .A1(n171), .B0(n168), .B1(IR[2]), .C0(
        muxres1[4]), .C1(n76), .Y(n81) );
  CLKINVX1 U393 ( .A(n82), .Y(n206) );
  AOI222XL U394 ( .A0(ReadData1[3]), .A1(n171), .B0(n75), .B1(IR[1]), .C0(
        muxres1[3]), .C1(n76), .Y(n82) );
  AOI221XL U395 ( .A0(n208), .A1(n173), .B0(RegDst[0]), .B1(IR[12]), .C0(
        RegDst[1]), .Y(n109) );
  AOI221XL U396 ( .A0(n208), .A1(n172), .B0(RegDst[0]), .B1(IR[11]), .C0(
        RegDst[1]), .Y(n110) );
  AOI221XL U397 ( .A0(n208), .A1(n174), .B0(RegDst[0]), .B1(IR[13]), .C0(
        RegDst[1]), .Y(n108) );
  NOR2BX1 U398 ( .AN(MemToReg[0]), .B(n170), .Y(n167) );
  NOR2BX1 U399 ( .AN(MemToReg[0]), .B(n170), .Y(n166) );
  NOR2BX1 U400 ( .AN(Jump), .B(n171), .Y(n75) );
  NOR2BX1 U401 ( .AN(Jump), .B(n171), .Y(n168) );
  NOR2BX1 U402 ( .AN(Jump), .B(n171), .Y(n169) );
  NOR2BX1 U403 ( .AN(MemToReg[0]), .B(n170), .Y(n113) );
  CLKBUFX3 U404 ( .A(rst_n), .Y(n179) );
  CLKINVX1 U405 ( .A(n106), .Y(n67) );
  AOI221XL U406 ( .A0(n208), .A1(IR[20]), .B0(RegDst[0]), .B1(IR[15]), .C0(
        RegDst[1]), .Y(n106) );
  CLKBUFX3 U407 ( .A(Jr), .Y(n171) );
  CLKINVX1 U408 ( .A(n107), .Y(n68) );
  AOI221XL U409 ( .A0(n208), .A1(n175), .B0(RegDst[0]), .B1(IR[14]), .C0(
        RegDst[1]), .Y(n107) );
  CLKBUFX3 U410 ( .A(MemToReg[1]), .Y(n170) );
  NOR2X1 U411 ( .A(MemRead), .B(MemWrite), .Y(CEN) );
  CLKBUFX3 U412 ( .A(IR[19]), .Y(n175) );
  CLKBUFX3 U413 ( .A(IR[18]), .Y(n174) );
  CLKBUFX3 U414 ( .A(IR[24]), .Y(n178) );
  CLKINVX1 U415 ( .A(RegDst[0]), .Y(n208) );
  CLKBUFX3 U416 ( .A(IR[16]), .Y(n172) );
  CLKBUFX3 U417 ( .A(IR[21]), .Y(n176) );
  CLKBUFX3 U418 ( .A(IR[17]), .Y(n173) );
  CLKBUFX3 U419 ( .A(IR[22]), .Y(n177) );
  NOR2BX1 U420 ( .AN(IR[8]), .B(n160), .Y(N36) );
  NOR2BX1 U421 ( .AN(IR[9]), .B(n161), .Y(N37) );
  NOR2BX1 U422 ( .AN(IR[10]), .B(n160), .Y(N38) );
  NOR2BX1 U423 ( .AN(IR[11]), .B(n161), .Y(N39) );
  NOR2BX1 U424 ( .AN(IR[12]), .B(n160), .Y(N40) );
  NOR2BX1 U425 ( .AN(IR[13]), .B(n161), .Y(N41) );
  NOR2BX1 U426 ( .AN(IR[14]), .B(n161), .Y(N42) );
  NOR2BX1 U427 ( .AN(IR[0]), .B(n162), .Y(N28) );
  NOR2BX1 U428 ( .AN(IR[1]), .B(n162), .Y(N29) );
  NOR2BX1 U429 ( .AN(IR[2]), .B(n160), .Y(N30) );
  NOR2BX1 U430 ( .AN(IR[3]), .B(n161), .Y(N31) );
  NOR2BX1 U431 ( .AN(IR[4]), .B(n160), .Y(N32) );
  NOR2BX1 U432 ( .AN(IR[5]), .B(n161), .Y(N33) );
  NOR2BX1 U433 ( .AN(IR[6]), .B(n160), .Y(N34) );
  NOR2BX1 U434 ( .AN(IR[7]), .B(n161), .Y(N35) );
endmodule

