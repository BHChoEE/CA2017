
module cache ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N42, N43, N44, N45, N46, \block[7][3][31] , \block[7][3][30] ,
         \block[7][3][29] , \block[7][3][28] , \block[7][3][27] ,
         \block[7][3][26] , \block[7][3][25] , \block[7][3][24] ,
         \block[7][3][23] , \block[7][3][22] , \block[7][3][21] ,
         \block[7][3][20] , \block[7][3][19] , \block[7][3][18] ,
         \block[7][3][17] , \block[7][3][16] , \block[7][3][15] ,
         \block[7][3][14] , \block[7][3][13] , \block[7][3][12] ,
         \block[7][3][11] , \block[7][3][10] , \block[7][3][9] ,
         \block[7][3][8] , \block[7][3][7] , \block[7][3][6] ,
         \block[7][3][5] , \block[7][3][4] , \block[7][3][3] ,
         \block[7][3][2] , \block[7][3][1] , \block[7][3][0] ,
         \block[7][2][31] , \block[7][2][30] , \block[7][2][29] ,
         \block[7][2][28] , \block[7][2][27] , \block[7][2][26] ,
         \block[7][2][25] , \block[7][2][24] , \block[7][2][23] ,
         \block[7][2][22] , \block[7][2][21] , \block[7][2][20] ,
         \block[7][2][19] , \block[7][2][18] , \block[7][2][17] ,
         \block[7][2][16] , \block[7][2][15] , \block[7][2][14] ,
         \block[7][2][13] , \block[7][2][12] , \block[7][2][11] ,
         \block[7][2][10] , \block[7][2][9] , \block[7][2][8] ,
         \block[7][2][7] , \block[7][2][6] , \block[7][2][5] ,
         \block[7][2][4] , \block[7][2][3] , \block[7][2][2] ,
         \block[7][2][1] , \block[7][2][0] , \block[7][1][31] ,
         \block[7][1][30] , \block[7][1][29] , \block[7][1][28] ,
         \block[7][1][27] , \block[7][1][26] , \block[7][1][25] ,
         \block[7][1][24] , \block[7][1][23] , \block[7][1][22] ,
         \block[7][1][21] , \block[7][1][20] , \block[7][1][19] ,
         \block[7][1][18] , \block[7][1][17] , \block[7][1][16] ,
         \block[7][1][15] , \block[7][1][14] , \block[7][1][13] ,
         \block[7][1][12] , \block[7][1][11] , \block[7][1][10] ,
         \block[7][1][9] , \block[7][1][8] , \block[7][1][7] ,
         \block[7][1][6] , \block[7][1][5] , \block[7][1][4] ,
         \block[7][1][3] , \block[7][1][2] , \block[7][1][1] ,
         \block[7][1][0] , \block[7][0][31] , \block[7][0][30] ,
         \block[7][0][29] , \block[7][0][28] , \block[7][0][27] ,
         \block[7][0][26] , \block[7][0][25] , \block[7][0][24] ,
         \block[7][0][23] , \block[7][0][22] , \block[7][0][21] ,
         \block[7][0][20] , \block[7][0][19] , \block[7][0][18] ,
         \block[7][0][17] , \block[7][0][16] , \block[7][0][15] ,
         \block[7][0][14] , \block[7][0][13] , \block[7][0][12] ,
         \block[7][0][11] , \block[7][0][10] , \block[7][0][9] ,
         \block[7][0][8] , \block[7][0][7] , \block[7][0][6] ,
         \block[7][0][5] , \block[7][0][4] , \block[7][0][3] ,
         \block[7][0][2] , \block[7][0][1] , \block[7][0][0] ,
         \block[6][3][31] , \block[6][3][30] , \block[6][3][29] ,
         \block[6][3][28] , \block[6][3][27] , \block[6][3][26] ,
         \block[6][3][25] , \block[6][3][24] , \block[6][3][23] ,
         \block[6][3][22] , \block[6][3][21] , \block[6][3][20] ,
         \block[6][3][19] , \block[6][3][18] , \block[6][3][17] ,
         \block[6][3][16] , \block[6][3][15] , \block[6][3][14] ,
         \block[6][3][13] , \block[6][3][12] , \block[6][3][11] ,
         \block[6][3][10] , \block[6][3][9] , \block[6][3][8] ,
         \block[6][3][7] , \block[6][3][6] , \block[6][3][5] ,
         \block[6][3][4] , \block[6][3][3] , \block[6][3][2] ,
         \block[6][3][1] , \block[6][3][0] , \block[6][2][31] ,
         \block[6][2][30] , \block[6][2][29] , \block[6][2][28] ,
         \block[6][2][27] , \block[6][2][26] , \block[6][2][25] ,
         \block[6][2][24] , \block[6][2][23] , \block[6][2][22] ,
         \block[6][2][21] , \block[6][2][20] , \block[6][2][19] ,
         \block[6][2][18] , \block[6][2][17] , \block[6][2][16] ,
         \block[6][2][15] , \block[6][2][14] , \block[6][2][13] ,
         \block[6][2][12] , \block[6][2][11] , \block[6][2][10] ,
         \block[6][2][9] , \block[6][2][8] , \block[6][2][7] ,
         \block[6][2][6] , \block[6][2][5] , \block[6][2][4] ,
         \block[6][2][3] , \block[6][2][2] , \block[6][2][1] ,
         \block[6][2][0] , \block[6][1][31] , \block[6][1][30] ,
         \block[6][1][29] , \block[6][1][28] , \block[6][1][27] ,
         \block[6][1][26] , \block[6][1][25] , \block[6][1][24] ,
         \block[6][1][23] , \block[6][1][22] , \block[6][1][21] ,
         \block[6][1][20] , \block[6][1][19] , \block[6][1][18] ,
         \block[6][1][17] , \block[6][1][16] , \block[6][1][15] ,
         \block[6][1][14] , \block[6][1][13] , \block[6][1][12] ,
         \block[6][1][11] , \block[6][1][10] , \block[6][1][9] ,
         \block[6][1][8] , \block[6][1][7] , \block[6][1][6] ,
         \block[6][1][5] , \block[6][1][4] , \block[6][1][3] ,
         \block[6][1][2] , \block[6][1][1] , \block[6][1][0] ,
         \block[6][0][31] , \block[6][0][30] , \block[6][0][29] ,
         \block[6][0][28] , \block[6][0][27] , \block[6][0][26] ,
         \block[6][0][25] , \block[6][0][24] , \block[6][0][23] ,
         \block[6][0][22] , \block[6][0][21] , \block[6][0][20] ,
         \block[6][0][19] , \block[6][0][18] , \block[6][0][17] ,
         \block[6][0][16] , \block[6][0][15] , \block[6][0][14] ,
         \block[6][0][13] , \block[6][0][12] , \block[6][0][11] ,
         \block[6][0][10] , \block[6][0][9] , \block[6][0][8] ,
         \block[6][0][7] , \block[6][0][6] , \block[6][0][5] ,
         \block[6][0][4] , \block[6][0][3] , \block[6][0][2] ,
         \block[6][0][1] , \block[6][0][0] , \block[5][3][31] ,
         \block[5][3][30] , \block[5][3][29] , \block[5][3][28] ,
         \block[5][3][27] , \block[5][3][26] , \block[5][3][25] ,
         \block[5][3][24] , \block[5][3][23] , \block[5][3][22] ,
         \block[5][3][21] , \block[5][3][20] , \block[5][3][19] ,
         \block[5][3][18] , \block[5][3][17] , \block[5][3][16] ,
         \block[5][3][15] , \block[5][3][14] , \block[5][3][13] ,
         \block[5][3][12] , \block[5][3][11] , \block[5][3][10] ,
         \block[5][3][9] , \block[5][3][8] , \block[5][3][7] ,
         \block[5][3][6] , \block[5][3][5] , \block[5][3][4] ,
         \block[5][3][3] , \block[5][3][2] , \block[5][3][1] ,
         \block[5][3][0] , \block[5][2][31] , \block[5][2][30] ,
         \block[5][2][29] , \block[5][2][28] , \block[5][2][27] ,
         \block[5][2][26] , \block[5][2][25] , \block[5][2][24] ,
         \block[5][2][23] , \block[5][2][22] , \block[5][2][21] ,
         \block[5][2][20] , \block[5][2][19] , \block[5][2][18] ,
         \block[5][2][17] , \block[5][2][16] , \block[5][2][15] ,
         \block[5][2][14] , \block[5][2][13] , \block[5][2][12] ,
         \block[5][2][11] , \block[5][2][10] , \block[5][2][9] ,
         \block[5][2][8] , \block[5][2][7] , \block[5][2][6] ,
         \block[5][2][5] , \block[5][2][4] , \block[5][2][3] ,
         \block[5][2][2] , \block[5][2][1] , \block[5][2][0] ,
         \block[5][1][31] , \block[5][1][30] , \block[5][1][29] ,
         \block[5][1][28] , \block[5][1][27] , \block[5][1][26] ,
         \block[5][1][25] , \block[5][1][24] , \block[5][1][23] ,
         \block[5][1][22] , \block[5][1][21] , \block[5][1][20] ,
         \block[5][1][19] , \block[5][1][18] , \block[5][1][17] ,
         \block[5][1][16] , \block[5][1][15] , \block[5][1][14] ,
         \block[5][1][13] , \block[5][1][12] , \block[5][1][11] ,
         \block[5][1][10] , \block[5][1][9] , \block[5][1][8] ,
         \block[5][1][7] , \block[5][1][6] , \block[5][1][5] ,
         \block[5][1][4] , \block[5][1][3] , \block[5][1][2] ,
         \block[5][1][1] , \block[5][1][0] , \block[5][0][31] ,
         \block[5][0][30] , \block[5][0][29] , \block[5][0][28] ,
         \block[5][0][27] , \block[5][0][26] , \block[5][0][25] ,
         \block[5][0][24] , \block[5][0][23] , \block[5][0][22] ,
         \block[5][0][21] , \block[5][0][20] , \block[5][0][19] ,
         \block[5][0][18] , \block[5][0][17] , \block[5][0][16] ,
         \block[5][0][15] , \block[5][0][14] , \block[5][0][13] ,
         \block[5][0][12] , \block[5][0][11] , \block[5][0][10] ,
         \block[5][0][9] , \block[5][0][8] , \block[5][0][7] ,
         \block[5][0][6] , \block[5][0][5] , \block[5][0][4] ,
         \block[5][0][3] , \block[5][0][2] , \block[5][0][1] ,
         \block[5][0][0] , \block[4][3][31] , \block[4][3][30] ,
         \block[4][3][29] , \block[4][3][28] , \block[4][3][27] ,
         \block[4][3][26] , \block[4][3][25] , \block[4][3][24] ,
         \block[4][3][23] , \block[4][3][22] , \block[4][3][21] ,
         \block[4][3][20] , \block[4][3][19] , \block[4][3][18] ,
         \block[4][3][17] , \block[4][3][16] , \block[4][3][15] ,
         \block[4][3][14] , \block[4][3][13] , \block[4][3][12] ,
         \block[4][3][11] , \block[4][3][10] , \block[4][3][9] ,
         \block[4][3][8] , \block[4][3][7] , \block[4][3][6] ,
         \block[4][3][5] , \block[4][3][4] , \block[4][3][3] ,
         \block[4][3][2] , \block[4][3][1] , \block[4][3][0] ,
         \block[4][2][31] , \block[4][2][30] , \block[4][2][29] ,
         \block[4][2][28] , \block[4][2][27] , \block[4][2][26] ,
         \block[4][2][25] , \block[4][2][24] , \block[4][2][23] ,
         \block[4][2][22] , \block[4][2][21] , \block[4][2][20] ,
         \block[4][2][19] , \block[4][2][18] , \block[4][2][17] ,
         \block[4][2][16] , \block[4][2][15] , \block[4][2][14] ,
         \block[4][2][13] , \block[4][2][12] , \block[4][2][11] ,
         \block[4][2][10] , \block[4][2][9] , \block[4][2][8] ,
         \block[4][2][7] , \block[4][2][6] , \block[4][2][5] ,
         \block[4][2][4] , \block[4][2][3] , \block[4][2][2] ,
         \block[4][2][1] , \block[4][2][0] , \block[4][1][31] ,
         \block[4][1][30] , \block[4][1][29] , \block[4][1][28] ,
         \block[4][1][27] , \block[4][1][26] , \block[4][1][25] ,
         \block[4][1][24] , \block[4][1][23] , \block[4][1][22] ,
         \block[4][1][21] , \block[4][1][20] , \block[4][1][19] ,
         \block[4][1][18] , \block[4][1][17] , \block[4][1][16] ,
         \block[4][1][15] , \block[4][1][14] , \block[4][1][13] ,
         \block[4][1][12] , \block[4][1][11] , \block[4][1][10] ,
         \block[4][1][9] , \block[4][1][8] , \block[4][1][7] ,
         \block[4][1][6] , \block[4][1][5] , \block[4][1][4] ,
         \block[4][1][3] , \block[4][1][2] , \block[4][1][1] ,
         \block[4][1][0] , \block[4][0][31] , \block[4][0][30] ,
         \block[4][0][29] , \block[4][0][28] , \block[4][0][27] ,
         \block[4][0][26] , \block[4][0][25] , \block[4][0][24] ,
         \block[4][0][23] , \block[4][0][22] , \block[4][0][21] ,
         \block[4][0][20] , \block[4][0][19] , \block[4][0][18] ,
         \block[4][0][17] , \block[4][0][16] , \block[4][0][15] ,
         \block[4][0][14] , \block[4][0][13] , \block[4][0][12] ,
         \block[4][0][11] , \block[4][0][10] , \block[4][0][9] ,
         \block[4][0][8] , \block[4][0][7] , \block[4][0][6] ,
         \block[4][0][5] , \block[4][0][4] , \block[4][0][3] ,
         \block[4][0][2] , \block[4][0][1] , \block[4][0][0] ,
         \block[3][3][31] , \block[3][3][30] , \block[3][3][29] ,
         \block[3][3][28] , \block[3][3][27] , \block[3][3][26] ,
         \block[3][3][25] , \block[3][3][24] , \block[3][3][23] ,
         \block[3][3][22] , \block[3][3][21] , \block[3][3][20] ,
         \block[3][3][19] , \block[3][3][18] , \block[3][3][17] ,
         \block[3][3][16] , \block[3][3][15] , \block[3][3][14] ,
         \block[3][3][13] , \block[3][3][12] , \block[3][3][11] ,
         \block[3][3][10] , \block[3][3][9] , \block[3][3][8] ,
         \block[3][3][7] , \block[3][3][6] , \block[3][3][5] ,
         \block[3][3][4] , \block[3][3][3] , \block[3][3][2] ,
         \block[3][3][1] , \block[3][3][0] , \block[3][2][31] ,
         \block[3][2][30] , \block[3][2][29] , \block[3][2][28] ,
         \block[3][2][27] , \block[3][2][26] , \block[3][2][25] ,
         \block[3][2][24] , \block[3][2][23] , \block[3][2][22] ,
         \block[3][2][21] , \block[3][2][20] , \block[3][2][19] ,
         \block[3][2][18] , \block[3][2][17] , \block[3][2][16] ,
         \block[3][2][15] , \block[3][2][14] , \block[3][2][13] ,
         \block[3][2][12] , \block[3][2][11] , \block[3][2][10] ,
         \block[3][2][9] , \block[3][2][8] , \block[3][2][7] ,
         \block[3][2][6] , \block[3][2][5] , \block[3][2][4] ,
         \block[3][2][3] , \block[3][2][2] , \block[3][2][1] ,
         \block[3][2][0] , \block[3][1][31] , \block[3][1][30] ,
         \block[3][1][29] , \block[3][1][28] , \block[3][1][27] ,
         \block[3][1][26] , \block[3][1][25] , \block[3][1][24] ,
         \block[3][1][23] , \block[3][1][22] , \block[3][1][21] ,
         \block[3][1][20] , \block[3][1][19] , \block[3][1][18] ,
         \block[3][1][17] , \block[3][1][16] , \block[3][1][15] ,
         \block[3][1][14] , \block[3][1][13] , \block[3][1][12] ,
         \block[3][1][11] , \block[3][1][10] , \block[3][1][9] ,
         \block[3][1][8] , \block[3][1][7] , \block[3][1][6] ,
         \block[3][1][5] , \block[3][1][4] , \block[3][1][3] ,
         \block[3][1][2] , \block[3][1][1] , \block[3][1][0] ,
         \block[3][0][31] , \block[3][0][30] , \block[3][0][29] ,
         \block[3][0][28] , \block[3][0][27] , \block[3][0][26] ,
         \block[3][0][25] , \block[3][0][24] , \block[3][0][23] ,
         \block[3][0][22] , \block[3][0][21] , \block[3][0][20] ,
         \block[3][0][19] , \block[3][0][18] , \block[3][0][17] ,
         \block[3][0][16] , \block[3][0][15] , \block[3][0][14] ,
         \block[3][0][13] , \block[3][0][12] , \block[3][0][11] ,
         \block[3][0][10] , \block[3][0][9] , \block[3][0][8] ,
         \block[3][0][7] , \block[3][0][6] , \block[3][0][5] ,
         \block[3][0][4] , \block[3][0][3] , \block[3][0][2] ,
         \block[3][0][1] , \block[3][0][0] , \block[2][3][31] ,
         \block[2][3][30] , \block[2][3][29] , \block[2][3][28] ,
         \block[2][3][27] , \block[2][3][26] , \block[2][3][25] ,
         \block[2][3][24] , \block[2][3][23] , \block[2][3][22] ,
         \block[2][3][21] , \block[2][3][20] , \block[2][3][19] ,
         \block[2][3][18] , \block[2][3][17] , \block[2][3][16] ,
         \block[2][3][15] , \block[2][3][14] , \block[2][3][13] ,
         \block[2][3][12] , \block[2][3][11] , \block[2][3][10] ,
         \block[2][3][9] , \block[2][3][8] , \block[2][3][7] ,
         \block[2][3][6] , \block[2][3][5] , \block[2][3][4] ,
         \block[2][3][3] , \block[2][3][2] , \block[2][3][1] ,
         \block[2][3][0] , \block[2][2][31] , \block[2][2][30] ,
         \block[2][2][29] , \block[2][2][28] , \block[2][2][27] ,
         \block[2][2][26] , \block[2][2][25] , \block[2][2][24] ,
         \block[2][2][23] , \block[2][2][22] , \block[2][2][21] ,
         \block[2][2][20] , \block[2][2][19] , \block[2][2][18] ,
         \block[2][2][17] , \block[2][2][16] , \block[2][2][15] ,
         \block[2][2][14] , \block[2][2][13] , \block[2][2][12] ,
         \block[2][2][11] , \block[2][2][10] , \block[2][2][9] ,
         \block[2][2][8] , \block[2][2][7] , \block[2][2][6] ,
         \block[2][2][5] , \block[2][2][4] , \block[2][2][3] ,
         \block[2][2][2] , \block[2][2][1] , \block[2][2][0] ,
         \block[2][1][31] , \block[2][1][30] , \block[2][1][29] ,
         \block[2][1][28] , \block[2][1][27] , \block[2][1][26] ,
         \block[2][1][25] , \block[2][1][24] , \block[2][1][23] ,
         \block[2][1][22] , \block[2][1][21] , \block[2][1][20] ,
         \block[2][1][19] , \block[2][1][18] , \block[2][1][17] ,
         \block[2][1][16] , \block[2][1][15] , \block[2][1][14] ,
         \block[2][1][13] , \block[2][1][12] , \block[2][1][11] ,
         \block[2][1][10] , \block[2][1][9] , \block[2][1][8] ,
         \block[2][1][7] , \block[2][1][6] , \block[2][1][5] ,
         \block[2][1][4] , \block[2][1][3] , \block[2][1][2] ,
         \block[2][1][1] , \block[2][1][0] , \block[2][0][31] ,
         \block[2][0][30] , \block[2][0][29] , \block[2][0][28] ,
         \block[2][0][27] , \block[2][0][26] , \block[2][0][25] ,
         \block[2][0][24] , \block[2][0][23] , \block[2][0][22] ,
         \block[2][0][21] , \block[2][0][20] , \block[2][0][19] ,
         \block[2][0][18] , \block[2][0][17] , \block[2][0][16] ,
         \block[2][0][15] , \block[2][0][14] , \block[2][0][13] ,
         \block[2][0][12] , \block[2][0][11] , \block[2][0][10] ,
         \block[2][0][9] , \block[2][0][8] , \block[2][0][7] ,
         \block[2][0][6] , \block[2][0][5] , \block[2][0][4] ,
         \block[2][0][3] , \block[2][0][2] , \block[2][0][1] ,
         \block[2][0][0] , \block[1][3][31] , \block[1][3][30] ,
         \block[1][3][29] , \block[1][3][28] , \block[1][3][27] ,
         \block[1][3][26] , \block[1][3][25] , \block[1][3][24] ,
         \block[1][3][23] , \block[1][3][22] , \block[1][3][21] ,
         \block[1][3][20] , \block[1][3][19] , \block[1][3][18] ,
         \block[1][3][17] , \block[1][3][16] , \block[1][3][15] ,
         \block[1][3][14] , \block[1][3][13] , \block[1][3][12] ,
         \block[1][3][11] , \block[1][3][10] , \block[1][3][9] ,
         \block[1][3][8] , \block[1][3][7] , \block[1][3][6] ,
         \block[1][3][5] , \block[1][3][4] , \block[1][3][3] ,
         \block[1][3][2] , \block[1][3][1] , \block[1][3][0] ,
         \block[1][2][31] , \block[1][2][30] , \block[1][2][29] ,
         \block[1][2][28] , \block[1][2][27] , \block[1][2][26] ,
         \block[1][2][25] , \block[1][2][24] , \block[1][2][23] ,
         \block[1][2][22] , \block[1][2][21] , \block[1][2][20] ,
         \block[1][2][19] , \block[1][2][18] , \block[1][2][17] ,
         \block[1][2][16] , \block[1][2][15] , \block[1][2][14] ,
         \block[1][2][13] , \block[1][2][12] , \block[1][2][11] ,
         \block[1][2][10] , \block[1][2][9] , \block[1][2][8] ,
         \block[1][2][7] , \block[1][2][6] , \block[1][2][5] ,
         \block[1][2][4] , \block[1][2][3] , \block[1][2][2] ,
         \block[1][2][1] , \block[1][2][0] , \block[1][1][31] ,
         \block[1][1][30] , \block[1][1][29] , \block[1][1][28] ,
         \block[1][1][27] , \block[1][1][26] , \block[1][1][25] ,
         \block[1][1][24] , \block[1][1][23] , \block[1][1][22] ,
         \block[1][1][21] , \block[1][1][20] , \block[1][1][19] ,
         \block[1][1][18] , \block[1][1][17] , \block[1][1][16] ,
         \block[1][1][15] , \block[1][1][14] , \block[1][1][13] ,
         \block[1][1][12] , \block[1][1][11] , \block[1][1][10] ,
         \block[1][1][9] , \block[1][1][8] , \block[1][1][7] ,
         \block[1][1][6] , \block[1][1][5] , \block[1][1][4] ,
         \block[1][1][3] , \block[1][1][2] , \block[1][1][1] ,
         \block[1][1][0] , \block[1][0][31] , \block[1][0][30] ,
         \block[1][0][29] , \block[1][0][28] , \block[1][0][27] ,
         \block[1][0][26] , \block[1][0][25] , \block[1][0][24] ,
         \block[1][0][23] , \block[1][0][22] , \block[1][0][21] ,
         \block[1][0][20] , \block[1][0][19] , \block[1][0][18] ,
         \block[1][0][17] , \block[1][0][16] , \block[1][0][15] ,
         \block[1][0][14] , \block[1][0][13] , \block[1][0][12] ,
         \block[1][0][11] , \block[1][0][10] , \block[1][0][9] ,
         \block[1][0][8] , \block[1][0][7] , \block[1][0][6] ,
         \block[1][0][5] , \block[1][0][4] , \block[1][0][3] ,
         \block[1][0][2] , \block[1][0][1] , \block[1][0][0] ,
         \block[0][3][31] , \block[0][3][30] , \block[0][3][29] ,
         \block[0][3][28] , \block[0][3][27] , \block[0][3][26] ,
         \block[0][3][25] , \block[0][3][24] , \block[0][3][23] ,
         \block[0][3][22] , \block[0][3][21] , \block[0][3][20] ,
         \block[0][3][19] , \block[0][3][18] , \block[0][3][17] ,
         \block[0][3][16] , \block[0][3][15] , \block[0][3][14] ,
         \block[0][3][13] , \block[0][3][12] , \block[0][3][11] ,
         \block[0][3][10] , \block[0][3][9] , \block[0][3][8] ,
         \block[0][3][7] , \block[0][3][6] , \block[0][3][5] ,
         \block[0][3][4] , \block[0][3][3] , \block[0][3][2] ,
         \block[0][3][1] , \block[0][3][0] , \block[0][2][31] ,
         \block[0][2][30] , \block[0][2][29] , \block[0][2][28] ,
         \block[0][2][27] , \block[0][2][26] , \block[0][2][25] ,
         \block[0][2][24] , \block[0][2][23] , \block[0][2][22] ,
         \block[0][2][21] , \block[0][2][20] , \block[0][2][19] ,
         \block[0][2][18] , \block[0][2][17] , \block[0][2][16] ,
         \block[0][2][15] , \block[0][2][14] , \block[0][2][13] ,
         \block[0][2][12] , \block[0][2][11] , \block[0][2][10] ,
         \block[0][2][9] , \block[0][2][8] , \block[0][2][7] ,
         \block[0][2][6] , \block[0][2][5] , \block[0][2][4] ,
         \block[0][2][3] , \block[0][2][2] , \block[0][2][1] ,
         \block[0][2][0] , \block[0][1][31] , \block[0][1][30] ,
         \block[0][1][29] , \block[0][1][28] , \block[0][1][27] ,
         \block[0][1][26] , \block[0][1][25] , \block[0][1][24] ,
         \block[0][1][23] , \block[0][1][22] , \block[0][1][21] ,
         \block[0][1][20] , \block[0][1][19] , \block[0][1][18] ,
         \block[0][1][17] , \block[0][1][16] , \block[0][1][15] ,
         \block[0][1][14] , \block[0][1][13] , \block[0][1][12] ,
         \block[0][1][11] , \block[0][1][10] , \block[0][1][9] ,
         \block[0][1][8] , \block[0][1][7] , \block[0][1][6] ,
         \block[0][1][5] , \block[0][1][4] , \block[0][1][3] ,
         \block[0][1][2] , \block[0][1][1] , \block[0][1][0] ,
         \block[0][0][31] , \block[0][0][30] , \block[0][0][29] ,
         \block[0][0][28] , \block[0][0][27] , \block[0][0][26] ,
         \block[0][0][25] , \block[0][0][24] , \block[0][0][23] ,
         \block[0][0][22] , \block[0][0][21] , \block[0][0][20] ,
         \block[0][0][19] , \block[0][0][18] , \block[0][0][17] ,
         \block[0][0][16] , \block[0][0][15] , \block[0][0][14] ,
         \block[0][0][13] , \block[0][0][12] , \block[0][0][11] ,
         \block[0][0][10] , \block[0][0][9] , \block[0][0][8] ,
         \block[0][0][7] , \block[0][0][6] , \block[0][0][5] ,
         \block[0][0][4] , \block[0][0][3] , \block[0][0][2] ,
         \block[0][0][1] , \block[0][0][0] , N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         rw_status, \tag[7][24] , \tag[7][23] , \tag[7][22] , \tag[7][21] ,
         \tag[7][18] , \tag[7][16] , \tag[7][15] , \tag[7][14] , \tag[7][13] ,
         \tag[7][12] , \tag[7][11] , \tag[7][10] , \tag[7][9] , \tag[7][8] ,
         \tag[7][3] , \tag[7][1] , \tag[7][0] , \tag[6][24] , \tag[6][23] ,
         \tag[6][22] , \tag[6][21] , \tag[6][18] , \tag[6][16] , \tag[6][15] ,
         \tag[6][14] , \tag[6][13] , \tag[6][12] , \tag[6][11] , \tag[6][10] ,
         \tag[6][9] , \tag[6][8] , \tag[6][3] , \tag[6][1] , \tag[6][0] ,
         \tag[5][24] , \tag[5][23] , \tag[5][22] , \tag[5][21] , \tag[5][18] ,
         \tag[5][16] , \tag[5][15] , \tag[5][14] , \tag[5][13] , \tag[5][12] ,
         \tag[5][11] , \tag[5][10] , \tag[5][9] , \tag[5][8] , \tag[5][3] ,
         \tag[5][1] , \tag[5][0] , \tag[4][24] , \tag[4][23] , \tag[4][22] ,
         \tag[4][21] , \tag[4][18] , \tag[4][16] , \tag[4][15] , \tag[4][14] ,
         \tag[4][13] , \tag[4][12] , \tag[4][11] , \tag[4][10] , \tag[4][9] ,
         \tag[4][8] , \tag[4][3] , \tag[4][1] , \tag[4][0] , \tag[3][24] ,
         \tag[3][23] , \tag[3][22] , \tag[3][21] , \tag[3][18] , \tag[3][16] ,
         \tag[3][15] , \tag[3][14] , \tag[3][13] , \tag[3][12] , \tag[3][11] ,
         \tag[3][10] , \tag[3][9] , \tag[3][8] , \tag[3][3] , \tag[3][1] ,
         \tag[3][0] , \tag[2][24] , \tag[2][23] , \tag[2][22] , \tag[2][21] ,
         \tag[2][18] , \tag[2][16] , \tag[2][15] , \tag[2][14] , \tag[2][13] ,
         \tag[2][12] , \tag[2][11] , \tag[2][10] , \tag[2][9] , \tag[2][8] ,
         \tag[2][3] , \tag[2][1] , \tag[2][0] , \tag[1][24] , \tag[1][23] ,
         \tag[1][22] , \tag[1][21] , \tag[1][18] , \tag[1][16] , \tag[1][15] ,
         \tag[1][14] , \tag[1][13] , \tag[1][12] , \tag[1][11] , \tag[1][10] ,
         \tag[1][9] , \tag[1][8] , \tag[1][3] , \tag[1][1] , \tag[1][0] ,
         \tag[0][24] , \tag[0][23] , \tag[0][22] , \tag[0][21] , \tag[0][18] ,
         \tag[0][16] , \tag[0][15] , \tag[0][14] , \tag[0][13] , \tag[0][12] ,
         \tag[0][11] , \tag[0][10] , \tag[0][9] , \tag[0][8] , \tag[0][3] ,
         \tag[0][1] , \tag[0][0] , N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, n101, n102,
         n138, n139, n174, n184, n185, n190, n195, n197, n198, n199, n200,
         n202, n205, n208, n258, n260, n261, n265, n267, n268, n269, n270,
         n272, n274, n276, n278, n280, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n295, n297, n301, n302, n303, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307;
  wire   [7:0] valid;
  wire   [7:0] dirty;
  wire   [1:0] state;
  wire   [31:0] next_proc_wdata;
  assign N42 = proc_addr[2];
  assign N43 = proc_addr[3];
  assign N44 = proc_addr[4];
  assign N45 = proc_addr[0];
  assign N46 = proc_addr[1];

  DFFRX1 \prev_mem_addr_reg[27]  ( .D(n2813), .CK(clk), .RN(n3762), .Q(
        mem_addr[27]), .QN(n1350) );
  DFFRX1 \prev_mem_addr_reg[26]  ( .D(n2814), .CK(clk), .RN(n3762), .Q(
        mem_addr[26]), .QN(n1349) );
  DFFRX1 \prev_mem_addr_reg[25]  ( .D(n2815), .CK(clk), .RN(n3762), .Q(
        mem_addr[25]), .QN(n1348) );
  DFFRX1 \prev_mem_addr_reg[24]  ( .D(n2816), .CK(clk), .RN(n3762), .Q(
        mem_addr[24]), .QN(n1347) );
  DFFRX1 \prev_mem_addr_reg[23]  ( .D(n2817), .CK(clk), .RN(n3762), .Q(
        mem_addr[23]), .QN(n1346) );
  DFFRX1 \prev_mem_addr_reg[22]  ( .D(n2818), .CK(clk), .RN(n3762), .Q(
        mem_addr[22]), .QN(n1345) );
  DFFRX1 \prev_mem_addr_reg[21]  ( .D(n2819), .CK(clk), .RN(n3762), .Q(
        mem_addr[21]), .QN(n1344) );
  DFFRX1 \prev_mem_addr_reg[20]  ( .D(n2820), .CK(clk), .RN(n3762), .Q(
        mem_addr[20]), .QN(n1343) );
  DFFRX1 \prev_mem_addr_reg[19]  ( .D(n2821), .CK(clk), .RN(n3762), .Q(
        mem_addr[19]), .QN(n1342) );
  DFFRX1 \prev_mem_addr_reg[18]  ( .D(n2822), .CK(clk), .RN(n3762), .Q(
        mem_addr[18]), .QN(n1341) );
  DFFRX1 \prev_mem_addr_reg[17]  ( .D(n2823), .CK(clk), .RN(n3762), .Q(
        mem_addr[17]), .QN(n1340) );
  DFFRX1 \prev_mem_addr_reg[16]  ( .D(n2824), .CK(clk), .RN(n3762), .Q(
        mem_addr[16]), .QN(n1339) );
  DFFRX1 \prev_mem_addr_reg[15]  ( .D(n2825), .CK(clk), .RN(n3761), .Q(
        mem_addr[15]), .QN(n1338) );
  DFFRX1 \prev_mem_addr_reg[14]  ( .D(n2826), .CK(clk), .RN(n3761), .Q(
        mem_addr[14]), .QN(n1337) );
  DFFRX1 \prev_mem_addr_reg[13]  ( .D(n2827), .CK(clk), .RN(n3761), .Q(
        mem_addr[13]), .QN(n1336) );
  DFFRX1 \prev_mem_addr_reg[12]  ( .D(n2828), .CK(clk), .RN(n3761), .Q(
        mem_addr[12]), .QN(n1335) );
  DFFRX1 \prev_mem_addr_reg[11]  ( .D(n2829), .CK(clk), .RN(n3761), .Q(
        mem_addr[11]), .QN(n1334) );
  DFFRX1 \prev_mem_addr_reg[10]  ( .D(n2830), .CK(clk), .RN(n3761), .Q(
        mem_addr[10]), .QN(n1333) );
  DFFRX1 \prev_mem_addr_reg[9]  ( .D(n2831), .CK(clk), .RN(n3761), .Q(
        mem_addr[9]), .QN(n1332) );
  DFFRX1 \prev_mem_addr_reg[8]  ( .D(n2832), .CK(clk), .RN(n3761), .Q(
        mem_addr[8]), .QN(n1331) );
  DFFRX1 \prev_mem_addr_reg[7]  ( .D(n2833), .CK(clk), .RN(n3761), .Q(
        mem_addr[7]), .QN(n1330) );
  DFFRX1 \prev_mem_addr_reg[6]  ( .D(n2834), .CK(clk), .RN(n3761), .Q(
        mem_addr[6]), .QN(n1329) );
  DFFRX1 \prev_mem_addr_reg[5]  ( .D(n2835), .CK(clk), .RN(n3761), .Q(
        mem_addr[5]), .QN(n1328) );
  DFFRX1 \prev_mem_addr_reg[4]  ( .D(n2836), .CK(clk), .RN(n3761), .Q(
        mem_addr[4]), .QN(n1327) );
  DFFRX1 \prev_mem_addr_reg[3]  ( .D(n2837), .CK(clk), .RN(n3760), .Q(
        mem_addr[3]), .QN(n1326) );
  DFFRX1 \prev_mem_addr_reg[2]  ( .D(n2838), .CK(clk), .RN(n3760), .Q(
        mem_addr[2]), .QN(n1325) );
  DFFRX1 \prev_mem_addr_reg[1]  ( .D(n2839), .CK(clk), .RN(n3760), .Q(
        mem_addr[1]), .QN(n1324) );
  DFFRX1 \prev_mem_addr_reg[0]  ( .D(n2840), .CK(clk), .RN(n3760), .Q(
        mem_addr[0]), .QN(n1323) );
  DFFRX1 prev_mem_write_reg ( .D(n2969), .CK(clk), .RN(n3759), .Q(mem_write), 
        .QN(n1322) );
  DFFRX1 \prev_proc_rdata_reg[31]  ( .D(n2748), .CK(clk), .RN(n3673), .Q(
        proc_rdata[31]), .QN(n1382) );
  DFFRX1 \prev_proc_rdata_reg[30]  ( .D(n2749), .CK(clk), .RN(n3673), .Q(
        proc_rdata[30]), .QN(n1381) );
  DFFRX1 \prev_proc_rdata_reg[29]  ( .D(n2750), .CK(clk), .RN(n3673), .Q(
        proc_rdata[29]), .QN(n1380) );
  DFFRX1 \prev_proc_rdata_reg[28]  ( .D(n2751), .CK(clk), .RN(n3673), .Q(
        proc_rdata[28]), .QN(n1379) );
  DFFRX1 \prev_proc_rdata_reg[27]  ( .D(n2752), .CK(clk), .RN(n3673), .Q(
        proc_rdata[27]), .QN(n1378) );
  DFFRX1 \prev_proc_rdata_reg[26]  ( .D(n2753), .CK(clk), .RN(n3673), .Q(
        proc_rdata[26]), .QN(n1377) );
  DFFRX1 \prev_proc_rdata_reg[25]  ( .D(n2754), .CK(clk), .RN(n3673), .Q(
        proc_rdata[25]), .QN(n1376) );
  DFFRX1 \prev_proc_rdata_reg[24]  ( .D(n2755), .CK(clk), .RN(n3673), .Q(
        proc_rdata[24]), .QN(n1375) );
  DFFRX1 \prev_proc_rdata_reg[23]  ( .D(n2756), .CK(clk), .RN(n3673), .Q(
        proc_rdata[23]), .QN(n1374) );
  DFFRX1 \prev_proc_rdata_reg[22]  ( .D(n2757), .CK(clk), .RN(n3673), .Q(
        proc_rdata[22]), .QN(n1373) );
  DFFRX1 \prev_proc_rdata_reg[21]  ( .D(n2758), .CK(clk), .RN(n3672), .Q(
        proc_rdata[21]), .QN(n1372) );
  DFFRX1 \prev_proc_rdata_reg[20]  ( .D(n2759), .CK(clk), .RN(n3672), .Q(
        proc_rdata[20]), .QN(n1371) );
  DFFRX1 \prev_proc_rdata_reg[19]  ( .D(n2760), .CK(clk), .RN(n3672), .Q(
        proc_rdata[19]), .QN(n1370) );
  DFFRX1 \prev_proc_rdata_reg[18]  ( .D(n2761), .CK(clk), .RN(n3672), .Q(
        proc_rdata[18]), .QN(n1369) );
  DFFRX1 \prev_proc_rdata_reg[17]  ( .D(n2762), .CK(clk), .RN(n3672), .Q(
        proc_rdata[17]), .QN(n1368) );
  DFFRX1 \prev_proc_rdata_reg[16]  ( .D(n2763), .CK(clk), .RN(n3672), .Q(
        proc_rdata[16]), .QN(n1367) );
  DFFRX1 \prev_proc_rdata_reg[15]  ( .D(n2764), .CK(clk), .RN(n3672), .Q(
        proc_rdata[15]), .QN(n1366) );
  DFFRX1 \prev_proc_rdata_reg[14]  ( .D(n2765), .CK(clk), .RN(n3672), .Q(
        proc_rdata[14]), .QN(n1365) );
  DFFRX1 \prev_proc_rdata_reg[13]  ( .D(n2766), .CK(clk), .RN(n3672), .Q(
        proc_rdata[13]), .QN(n1364) );
  DFFRX1 \prev_proc_rdata_reg[12]  ( .D(n2767), .CK(clk), .RN(n3672), .Q(
        proc_rdata[12]), .QN(n1363) );
  DFFRX1 \prev_proc_rdata_reg[11]  ( .D(n2768), .CK(clk), .RN(n3672), .Q(
        proc_rdata[11]), .QN(n1362) );
  DFFRX1 \prev_proc_rdata_reg[10]  ( .D(n2769), .CK(clk), .RN(n3672), .Q(
        proc_rdata[10]), .QN(n1361) );
  DFFRX1 \prev_proc_rdata_reg[9]  ( .D(n2770), .CK(clk), .RN(n3671), .Q(
        proc_rdata[9]), .QN(n1360) );
  DFFRX1 \prev_proc_rdata_reg[8]  ( .D(n2771), .CK(clk), .RN(n3671), .Q(
        proc_rdata[8]), .QN(n1359) );
  DFFRX1 \prev_proc_rdata_reg[7]  ( .D(n2772), .CK(clk), .RN(n3671), .Q(
        proc_rdata[7]), .QN(n1358) );
  DFFRX1 \prev_proc_rdata_reg[6]  ( .D(n2773), .CK(clk), .RN(n3671), .Q(
        proc_rdata[6]), .QN(n1357) );
  DFFRX1 \prev_proc_rdata_reg[5]  ( .D(n2774), .CK(clk), .RN(n3671), .Q(
        proc_rdata[5]), .QN(n1356) );
  DFFRX1 \prev_proc_rdata_reg[4]  ( .D(n2775), .CK(clk), .RN(n3671), .Q(
        proc_rdata[4]), .QN(n1355) );
  DFFRX1 \prev_proc_rdata_reg[3]  ( .D(n2776), .CK(clk), .RN(n3671), .Q(
        proc_rdata[3]), .QN(n1354) );
  DFFRX1 \prev_proc_rdata_reg[2]  ( .D(n2777), .CK(clk), .RN(n3671), .Q(
        proc_rdata[2]), .QN(n1353) );
  DFFRX1 \prev_proc_rdata_reg[1]  ( .D(n2778), .CK(clk), .RN(n3671), .Q(
        proc_rdata[1]), .QN(n1352) );
  DFFRX1 \prev_proc_rdata_reg[0]  ( .D(n2779), .CK(clk), .RN(n3671), .Q(
        proc_rdata[0]), .QN(n1351) );
  DFFRX1 prev_proc_stall_reg ( .D(n1715), .CK(clk), .RN(n3671), .Q(proc_stall), 
        .QN(n1120) );
  DFFRX1 prev_mem_read_reg ( .D(n1714), .CK(clk), .RN(n3671), .Q(mem_read), 
        .QN(n1121) );
  DFFRX1 \block_reg[7][0][31]  ( .D(n1820), .CK(clk), .RN(n3751), .Q(
        \block[7][0][31] ), .QN(n1015) );
  DFFRX1 \block_reg[7][0][30]  ( .D(n1821), .CK(clk), .RN(n3751), .Q(
        \block[7][0][30] ), .QN(n1014) );
  DFFRX1 \block_reg[7][0][29]  ( .D(n1822), .CK(clk), .RN(n3750), .Q(
        \block[7][0][29] ), .QN(n1013) );
  DFFRX1 \block_reg[7][0][28]  ( .D(n1823), .CK(clk), .RN(n3750), .Q(
        \block[7][0][28] ), .QN(n1012) );
  DFFRX1 \block_reg[7][0][27]  ( .D(n1824), .CK(clk), .RN(n3750), .Q(
        \block[7][0][27] ), .QN(n1011) );
  DFFRX1 \block_reg[7][0][26]  ( .D(n1825), .CK(clk), .RN(n3750), .Q(
        \block[7][0][26] ), .QN(n1010) );
  DFFRX1 \block_reg[7][0][25]  ( .D(n1826), .CK(clk), .RN(n3750), .Q(
        \block[7][0][25] ), .QN(n1009) );
  DFFRX1 \block_reg[7][0][24]  ( .D(n1827), .CK(clk), .RN(n3750), .Q(
        \block[7][0][24] ), .QN(n1008) );
  DFFRX1 \block_reg[7][0][23]  ( .D(n1828), .CK(clk), .RN(n3750), .Q(
        \block[7][0][23] ), .QN(n1007) );
  DFFRX1 \block_reg[7][0][22]  ( .D(n1829), .CK(clk), .RN(n3750), .Q(
        \block[7][0][22] ), .QN(n1006) );
  DFFRX1 \block_reg[7][0][21]  ( .D(n1830), .CK(clk), .RN(n3750), .Q(
        \block[7][0][21] ), .QN(n1005) );
  DFFRX1 \block_reg[7][0][20]  ( .D(n1831), .CK(clk), .RN(n3750), .Q(
        \block[7][0][20] ), .QN(n1004) );
  DFFRX1 \block_reg[7][0][19]  ( .D(n1832), .CK(clk), .RN(n3750), .Q(
        \block[7][0][19] ), .QN(n1003) );
  DFFRX1 \block_reg[7][0][18]  ( .D(n1833), .CK(clk), .RN(n3750), .Q(
        \block[7][0][18] ), .QN(n1002) );
  DFFRX1 \block_reg[7][0][17]  ( .D(n1834), .CK(clk), .RN(n3749), .Q(
        \block[7][0][17] ), .QN(n1001) );
  DFFRX1 \block_reg[7][0][16]  ( .D(n1835), .CK(clk), .RN(n3749), .Q(
        \block[7][0][16] ), .QN(n1000) );
  DFFRX1 \block_reg[7][0][15]  ( .D(n1836), .CK(clk), .RN(n3749), .Q(
        \block[7][0][15] ), .QN(n999) );
  DFFRX1 \block_reg[7][0][14]  ( .D(n1837), .CK(clk), .RN(n3749), .Q(
        \block[7][0][14] ), .QN(n998) );
  DFFRX1 \block_reg[7][0][13]  ( .D(n1838), .CK(clk), .RN(n3749), .Q(
        \block[7][0][13] ), .QN(n997) );
  DFFRX1 \block_reg[7][0][12]  ( .D(n1839), .CK(clk), .RN(n3749), .Q(
        \block[7][0][12] ), .QN(n996) );
  DFFRX1 \block_reg[7][0][11]  ( .D(n1840), .CK(clk), .RN(n3749), .Q(
        \block[7][0][11] ), .QN(n995) );
  DFFRX1 \block_reg[7][0][10]  ( .D(n1841), .CK(clk), .RN(n3749), .Q(
        \block[7][0][10] ), .QN(n994) );
  DFFRX1 \block_reg[7][0][9]  ( .D(n1842), .CK(clk), .RN(n3749), .Q(
        \block[7][0][9] ), .QN(n993) );
  DFFRX1 \block_reg[7][0][8]  ( .D(n1843), .CK(clk), .RN(n3749), .Q(
        \block[7][0][8] ), .QN(n992) );
  DFFRX1 \block_reg[7][0][7]  ( .D(n1844), .CK(clk), .RN(n3749), .Q(
        \block[7][0][7] ), .QN(n991) );
  DFFRX1 \block_reg[7][0][6]  ( .D(n1845), .CK(clk), .RN(n3749), .Q(
        \block[7][0][6] ), .QN(n990) );
  DFFRX1 \block_reg[7][0][5]  ( .D(n1846), .CK(clk), .RN(n3748), .Q(
        \block[7][0][5] ), .QN(n989) );
  DFFRX1 \block_reg[7][0][4]  ( .D(n1847), .CK(clk), .RN(n3748), .Q(
        \block[7][0][4] ), .QN(n988) );
  DFFRX1 \block_reg[7][0][3]  ( .D(n1848), .CK(clk), .RN(n3748), .Q(
        \block[7][0][3] ), .QN(n987) );
  DFFRX1 \block_reg[7][0][2]  ( .D(n1849), .CK(clk), .RN(n3748), .Q(
        \block[7][0][2] ), .QN(n986) );
  DFFRX1 \block_reg[7][0][1]  ( .D(n1850), .CK(clk), .RN(n3748), .Q(
        \block[7][0][1] ), .QN(n985) );
  DFFRX1 \block_reg[7][0][0]  ( .D(n1851), .CK(clk), .RN(n3748), .Q(
        \block[7][0][0] ), .QN(n984) );
  DFFRX1 \block_reg[3][0][31]  ( .D(n2332), .CK(clk), .RN(n3740), .Q(
        \block[3][0][31] ), .QN(n503) );
  DFFRX1 \block_reg[3][0][30]  ( .D(n2333), .CK(clk), .RN(n3740), .Q(
        \block[3][0][30] ), .QN(n502) );
  DFFRX1 \block_reg[3][0][29]  ( .D(n2334), .CK(clk), .RN(n3740), .Q(
        \block[3][0][29] ), .QN(n501) );
  DFFRX1 \block_reg[3][0][28]  ( .D(n2335), .CK(clk), .RN(n3740), .Q(
        \block[3][0][28] ), .QN(n500) );
  DFFRX1 \block_reg[3][0][27]  ( .D(n2336), .CK(clk), .RN(n3740), .Q(
        \block[3][0][27] ), .QN(n499) );
  DFFRX1 \block_reg[3][0][26]  ( .D(n2337), .CK(clk), .RN(n3740), .Q(
        \block[3][0][26] ), .QN(n498) );
  DFFRX1 \block_reg[3][0][25]  ( .D(n2338), .CK(clk), .RN(n3739), .Q(
        \block[3][0][25] ), .QN(n497) );
  DFFRX1 \block_reg[3][0][24]  ( .D(n2339), .CK(clk), .RN(n3739), .Q(
        \block[3][0][24] ), .QN(n496) );
  DFFRX1 \block_reg[3][0][23]  ( .D(n2340), .CK(clk), .RN(n3739), .Q(
        \block[3][0][23] ), .QN(n495) );
  DFFRX1 \block_reg[3][0][22]  ( .D(n2341), .CK(clk), .RN(n3739), .Q(
        \block[3][0][22] ), .QN(n494) );
  DFFRX1 \block_reg[3][0][21]  ( .D(n2342), .CK(clk), .RN(n3739), .Q(
        \block[3][0][21] ), .QN(n493) );
  DFFRX1 \block_reg[3][0][20]  ( .D(n2343), .CK(clk), .RN(n3739), .Q(
        \block[3][0][20] ), .QN(n492) );
  DFFRX1 \block_reg[3][0][19]  ( .D(n2344), .CK(clk), .RN(n3739), .Q(
        \block[3][0][19] ), .QN(n491) );
  DFFRX1 \block_reg[3][0][18]  ( .D(n2345), .CK(clk), .RN(n3739), .Q(
        \block[3][0][18] ), .QN(n490) );
  DFFRX1 \block_reg[3][0][17]  ( .D(n2346), .CK(clk), .RN(n3739), .Q(
        \block[3][0][17] ), .QN(n489) );
  DFFRX1 \block_reg[3][0][16]  ( .D(n2347), .CK(clk), .RN(n3739), .Q(
        \block[3][0][16] ), .QN(n488) );
  DFFRX1 \block_reg[3][0][15]  ( .D(n2348), .CK(clk), .RN(n3739), .Q(
        \block[3][0][15] ), .QN(n487) );
  DFFRX1 \block_reg[3][0][14]  ( .D(n2349), .CK(clk), .RN(n3739), .Q(
        \block[3][0][14] ), .QN(n486) );
  DFFRX1 \block_reg[3][0][13]  ( .D(n2350), .CK(clk), .RN(n3738), .Q(
        \block[3][0][13] ), .QN(n485) );
  DFFRX1 \block_reg[3][0][12]  ( .D(n2351), .CK(clk), .RN(n3738), .Q(
        \block[3][0][12] ), .QN(n484) );
  DFFRX1 \block_reg[3][0][11]  ( .D(n2352), .CK(clk), .RN(n3738), .Q(
        \block[3][0][11] ), .QN(n483) );
  DFFRX1 \block_reg[3][0][10]  ( .D(n2353), .CK(clk), .RN(n3738), .Q(
        \block[3][0][10] ), .QN(n482) );
  DFFRX1 \block_reg[3][0][9]  ( .D(n2354), .CK(clk), .RN(n3738), .Q(
        \block[3][0][9] ), .QN(n481) );
  DFFRX1 \block_reg[3][0][8]  ( .D(n2355), .CK(clk), .RN(n3738), .Q(
        \block[3][0][8] ), .QN(n480) );
  DFFRX1 \block_reg[3][0][7]  ( .D(n2356), .CK(clk), .RN(n3738), .Q(
        \block[3][0][7] ), .QN(n479) );
  DFFRX1 \block_reg[3][0][6]  ( .D(n2357), .CK(clk), .RN(n3738), .Q(
        \block[3][0][6] ), .QN(n478) );
  DFFRX1 \block_reg[3][0][5]  ( .D(n2358), .CK(clk), .RN(n3738), .Q(
        \block[3][0][5] ), .QN(n477) );
  DFFRX1 \block_reg[3][0][4]  ( .D(n2359), .CK(clk), .RN(n3738), .Q(
        \block[3][0][4] ), .QN(n476) );
  DFFRX1 \block_reg[3][0][3]  ( .D(n2360), .CK(clk), .RN(n3738), .Q(
        \block[3][0][3] ), .QN(n475) );
  DFFRX1 \block_reg[3][0][2]  ( .D(n2361), .CK(clk), .RN(n3738), .Q(
        \block[3][0][2] ), .QN(n474) );
  DFFRX1 \block_reg[3][0][1]  ( .D(n2362), .CK(clk), .RN(n3737), .Q(
        \block[3][0][1] ), .QN(n473) );
  DFFRX1 \block_reg[3][0][0]  ( .D(n2363), .CK(clk), .RN(n3737), .Q(
        \block[3][0][0] ), .QN(n472) );
  DFFRX1 \block_reg[7][3][31]  ( .D(n1724), .CK(clk), .RN(n3732), .Q(
        \block[7][3][31] ), .QN(n1111) );
  DFFRX1 \block_reg[7][3][30]  ( .D(n1725), .CK(clk), .RN(n3732), .Q(
        \block[7][3][30] ), .QN(n1110) );
  DFFRX1 \block_reg[7][3][29]  ( .D(n1726), .CK(clk), .RN(n3732), .Q(
        \block[7][3][29] ), .QN(n1109) );
  DFFRX1 \block_reg[7][3][28]  ( .D(n1727), .CK(clk), .RN(n3732), .Q(
        \block[7][3][28] ), .QN(n1108) );
  DFFRX1 \block_reg[7][3][27]  ( .D(n1728), .CK(clk), .RN(n3732), .Q(
        \block[7][3][27] ), .QN(n1107) );
  DFFRX1 \block_reg[7][3][26]  ( .D(n1729), .CK(clk), .RN(n3732), .Q(
        \block[7][3][26] ), .QN(n1106) );
  DFFRX1 \block_reg[7][3][25]  ( .D(n1730), .CK(clk), .RN(n3731), .Q(
        \block[7][3][25] ), .QN(n1105) );
  DFFRX1 \block_reg[7][3][24]  ( .D(n1731), .CK(clk), .RN(n3731), .Q(
        \block[7][3][24] ), .QN(n1104) );
  DFFRX1 \block_reg[7][3][23]  ( .D(n1732), .CK(clk), .RN(n3731), .Q(
        \block[7][3][23] ), .QN(n1103) );
  DFFRX1 \block_reg[7][3][22]  ( .D(n1733), .CK(clk), .RN(n3731), .Q(
        \block[7][3][22] ), .QN(n1102) );
  DFFRX1 \block_reg[7][3][21]  ( .D(n1734), .CK(clk), .RN(n3731), .Q(
        \block[7][3][21] ), .QN(n1101) );
  DFFRX1 \block_reg[7][3][20]  ( .D(n1735), .CK(clk), .RN(n3731), .Q(
        \block[7][3][20] ), .QN(n1100) );
  DFFRX1 \block_reg[7][3][19]  ( .D(n1736), .CK(clk), .RN(n3731), .Q(
        \block[7][3][19] ), .QN(n1099) );
  DFFRX1 \block_reg[7][3][18]  ( .D(n1737), .CK(clk), .RN(n3731), .Q(
        \block[7][3][18] ), .QN(n1098) );
  DFFRX1 \block_reg[7][3][17]  ( .D(n1738), .CK(clk), .RN(n3731), .Q(
        \block[7][3][17] ), .QN(n1097) );
  DFFRX1 \block_reg[7][3][16]  ( .D(n1739), .CK(clk), .RN(n3731), .Q(
        \block[7][3][16] ), .QN(n1096) );
  DFFRX1 \block_reg[7][3][15]  ( .D(n1740), .CK(clk), .RN(n3731), .Q(
        \block[7][3][15] ), .QN(n1095) );
  DFFRX1 \block_reg[7][3][14]  ( .D(n1741), .CK(clk), .RN(n3731), .Q(
        \block[7][3][14] ), .QN(n1094) );
  DFFRX1 \block_reg[7][3][13]  ( .D(n1742), .CK(clk), .RN(n3730), .Q(
        \block[7][3][13] ), .QN(n1093) );
  DFFRX1 \block_reg[7][3][12]  ( .D(n1743), .CK(clk), .RN(n3730), .Q(
        \block[7][3][12] ), .QN(n1092) );
  DFFRX1 \block_reg[7][3][11]  ( .D(n1744), .CK(clk), .RN(n3730), .Q(
        \block[7][3][11] ), .QN(n1091) );
  DFFRX1 \block_reg[7][3][10]  ( .D(n1745), .CK(clk), .RN(n3730), .Q(
        \block[7][3][10] ), .QN(n1090) );
  DFFRX1 \block_reg[7][3][9]  ( .D(n1746), .CK(clk), .RN(n3730), .Q(
        \block[7][3][9] ), .QN(n1089) );
  DFFRX1 \block_reg[7][3][8]  ( .D(n1747), .CK(clk), .RN(n3730), .Q(
        \block[7][3][8] ), .QN(n1088) );
  DFFRX1 \block_reg[7][3][7]  ( .D(n1748), .CK(clk), .RN(n3730), .Q(
        \block[7][3][7] ), .QN(n1087) );
  DFFRX1 \block_reg[7][3][6]  ( .D(n1749), .CK(clk), .RN(n3730), .Q(
        \block[7][3][6] ), .QN(n1086) );
  DFFRX1 \block_reg[7][3][5]  ( .D(n1750), .CK(clk), .RN(n3730), .Q(
        \block[7][3][5] ), .QN(n1085) );
  DFFRX1 \block_reg[7][3][4]  ( .D(n1751), .CK(clk), .RN(n3730), .Q(
        \block[7][3][4] ), .QN(n1084) );
  DFFRX1 \block_reg[7][3][3]  ( .D(n1752), .CK(clk), .RN(n3730), .Q(
        \block[7][3][3] ), .QN(n1083) );
  DFFRX1 \block_reg[7][3][2]  ( .D(n1753), .CK(clk), .RN(n3730), .Q(
        \block[7][3][2] ), .QN(n1082) );
  DFFRX1 \block_reg[7][3][1]  ( .D(n1754), .CK(clk), .RN(n3729), .Q(
        \block[7][3][1] ), .QN(n1081) );
  DFFRX1 \block_reg[7][3][0]  ( .D(n1755), .CK(clk), .RN(n3729), .Q(
        \block[7][3][0] ), .QN(n1080) );
  DFFRX1 \block_reg[3][3][31]  ( .D(n2236), .CK(clk), .RN(n3721), .Q(
        \block[3][3][31] ), .QN(n599) );
  DFFRX1 \block_reg[3][3][30]  ( .D(n2237), .CK(clk), .RN(n3721), .Q(
        \block[3][3][30] ), .QN(n598) );
  DFFRX1 \block_reg[3][3][29]  ( .D(n2238), .CK(clk), .RN(n3721), .Q(
        \block[3][3][29] ), .QN(n597) );
  DFFRX1 \block_reg[3][3][28]  ( .D(n2239), .CK(clk), .RN(n3721), .Q(
        \block[3][3][28] ), .QN(n596) );
  DFFRX1 \block_reg[3][3][27]  ( .D(n2240), .CK(clk), .RN(n3721), .Q(
        \block[3][3][27] ), .QN(n595) );
  DFFRX1 \block_reg[3][3][26]  ( .D(n2241), .CK(clk), .RN(n3721), .Q(
        \block[3][3][26] ), .QN(n594) );
  DFFRX1 \block_reg[3][3][25]  ( .D(n2242), .CK(clk), .RN(n3721), .Q(
        \block[3][3][25] ), .QN(n593) );
  DFFRX1 \block_reg[3][3][24]  ( .D(n2243), .CK(clk), .RN(n3721), .Q(
        \block[3][3][24] ), .QN(n592) );
  DFFRX1 \block_reg[3][3][23]  ( .D(n2244), .CK(clk), .RN(n3721), .Q(
        \block[3][3][23] ), .QN(n591) );
  DFFRX1 \block_reg[3][3][22]  ( .D(n2245), .CK(clk), .RN(n3721), .Q(
        \block[3][3][22] ), .QN(n590) );
  DFFRX1 \block_reg[3][3][21]  ( .D(n2246), .CK(clk), .RN(n3720), .Q(
        \block[3][3][21] ), .QN(n589) );
  DFFRX1 \block_reg[3][3][20]  ( .D(n2247), .CK(clk), .RN(n3720), .Q(
        \block[3][3][20] ), .QN(n588) );
  DFFRX1 \block_reg[3][3][19]  ( .D(n2248), .CK(clk), .RN(n3720), .Q(
        \block[3][3][19] ), .QN(n587) );
  DFFRX1 \block_reg[3][3][18]  ( .D(n2249), .CK(clk), .RN(n3720), .Q(
        \block[3][3][18] ), .QN(n586) );
  DFFRX1 \block_reg[3][3][17]  ( .D(n2250), .CK(clk), .RN(n3720), .Q(
        \block[3][3][17] ), .QN(n585) );
  DFFRX1 \block_reg[3][3][16]  ( .D(n2251), .CK(clk), .RN(n3720), .Q(
        \block[3][3][16] ), .QN(n584) );
  DFFRX1 \block_reg[3][3][15]  ( .D(n2252), .CK(clk), .RN(n3720), .Q(
        \block[3][3][15] ), .QN(n583) );
  DFFRX1 \block_reg[3][3][14]  ( .D(n2253), .CK(clk), .RN(n3720), .Q(
        \block[3][3][14] ), .QN(n582) );
  DFFRX1 \block_reg[3][3][13]  ( .D(n2254), .CK(clk), .RN(n3720), .Q(
        \block[3][3][13] ), .QN(n581) );
  DFFRX1 \block_reg[3][3][12]  ( .D(n2255), .CK(clk), .RN(n3720), .Q(
        \block[3][3][12] ), .QN(n580) );
  DFFRX1 \block_reg[3][3][11]  ( .D(n2256), .CK(clk), .RN(n3720), .Q(
        \block[3][3][11] ), .QN(n579) );
  DFFRX1 \block_reg[3][3][10]  ( .D(n2257), .CK(clk), .RN(n3720), .Q(
        \block[3][3][10] ), .QN(n578) );
  DFFRX1 \block_reg[3][3][9]  ( .D(n2258), .CK(clk), .RN(n3719), .Q(
        \block[3][3][9] ), .QN(n577) );
  DFFRX1 \block_reg[3][3][8]  ( .D(n2259), .CK(clk), .RN(n3719), .Q(
        \block[3][3][8] ), .QN(n576) );
  DFFRX1 \block_reg[3][3][7]  ( .D(n2260), .CK(clk), .RN(n3719), .Q(
        \block[3][3][7] ), .QN(n575) );
  DFFRX1 \block_reg[3][3][6]  ( .D(n2261), .CK(clk), .RN(n3719), .Q(
        \block[3][3][6] ), .QN(n574) );
  DFFRX1 \block_reg[3][3][5]  ( .D(n2262), .CK(clk), .RN(n3719), .Q(
        \block[3][3][5] ), .QN(n573) );
  DFFRX1 \block_reg[3][3][4]  ( .D(n2263), .CK(clk), .RN(n3719), .Q(
        \block[3][3][4] ), .QN(n572) );
  DFFRX1 \block_reg[3][3][3]  ( .D(n2264), .CK(clk), .RN(n3719), .Q(
        \block[3][3][3] ), .QN(n571) );
  DFFRX1 \block_reg[3][3][2]  ( .D(n2265), .CK(clk), .RN(n3719), .Q(
        \block[3][3][2] ), .QN(n570) );
  DFFRX1 \block_reg[3][3][1]  ( .D(n2266), .CK(clk), .RN(n3719), .Q(
        \block[3][3][1] ), .QN(n569) );
  DFFRX1 \block_reg[3][3][0]  ( .D(n2267), .CK(clk), .RN(n3719), .Q(
        \block[3][3][0] ), .QN(n568) );
  DFFRX1 \block_reg[7][2][31]  ( .D(n1756), .CK(clk), .RN(n3711), .Q(
        \block[7][2][31] ), .QN(n1079) );
  DFFRX1 \block_reg[7][2][30]  ( .D(n1757), .CK(clk), .RN(n3711), .Q(
        \block[7][2][30] ), .QN(n1078) );
  DFFRX1 \block_reg[7][2][29]  ( .D(n1758), .CK(clk), .RN(n3710), .Q(
        \block[7][2][29] ), .QN(n1077) );
  DFFRX1 \block_reg[7][2][28]  ( .D(n1759), .CK(clk), .RN(n3710), .Q(
        \block[7][2][28] ), .QN(n1076) );
  DFFRX1 \block_reg[7][2][27]  ( .D(n1760), .CK(clk), .RN(n3710), .Q(
        \block[7][2][27] ), .QN(n1075) );
  DFFRX1 \block_reg[7][2][26]  ( .D(n1761), .CK(clk), .RN(n3710), .Q(
        \block[7][2][26] ), .QN(n1074) );
  DFFRX1 \block_reg[7][2][25]  ( .D(n1762), .CK(clk), .RN(n3710), .Q(
        \block[7][2][25] ), .QN(n1073) );
  DFFRX1 \block_reg[7][2][24]  ( .D(n1763), .CK(clk), .RN(n3710), .Q(
        \block[7][2][24] ), .QN(n1072) );
  DFFRX1 \block_reg[7][2][23]  ( .D(n1764), .CK(clk), .RN(n3710), .Q(
        \block[7][2][23] ), .QN(n1071) );
  DFFRX1 \block_reg[7][2][22]  ( .D(n1765), .CK(clk), .RN(n3710), .Q(
        \block[7][2][22] ), .QN(n1070) );
  DFFRX1 \block_reg[7][2][21]  ( .D(n1766), .CK(clk), .RN(n3710), .Q(
        \block[7][2][21] ), .QN(n1069) );
  DFFRX1 \block_reg[7][2][20]  ( .D(n1767), .CK(clk), .RN(n3710), .Q(
        \block[7][2][20] ), .QN(n1068) );
  DFFRX1 \block_reg[7][2][19]  ( .D(n1768), .CK(clk), .RN(n3710), .Q(
        \block[7][2][19] ), .QN(n1067) );
  DFFRX1 \block_reg[7][2][18]  ( .D(n1769), .CK(clk), .RN(n3710), .Q(
        \block[7][2][18] ), .QN(n1066) );
  DFFRX1 \block_reg[7][2][17]  ( .D(n1770), .CK(clk), .RN(n3709), .Q(
        \block[7][2][17] ), .QN(n1065) );
  DFFRX1 \block_reg[7][2][16]  ( .D(n1771), .CK(clk), .RN(n3709), .Q(
        \block[7][2][16] ), .QN(n1064) );
  DFFRX1 \block_reg[7][2][15]  ( .D(n1772), .CK(clk), .RN(n3709), .Q(
        \block[7][2][15] ), .QN(n1063) );
  DFFRX1 \block_reg[7][2][14]  ( .D(n1773), .CK(clk), .RN(n3709), .Q(
        \block[7][2][14] ), .QN(n1062) );
  DFFRX1 \block_reg[7][2][13]  ( .D(n1774), .CK(clk), .RN(n3709), .Q(
        \block[7][2][13] ), .QN(n1061) );
  DFFRX1 \block_reg[7][2][12]  ( .D(n1775), .CK(clk), .RN(n3709), .Q(
        \block[7][2][12] ), .QN(n1060) );
  DFFRX1 \block_reg[7][2][11]  ( .D(n1776), .CK(clk), .RN(n3709), .Q(
        \block[7][2][11] ), .QN(n1059) );
  DFFRX1 \block_reg[7][2][10]  ( .D(n1777), .CK(clk), .RN(n3709), .Q(
        \block[7][2][10] ), .QN(n1058) );
  DFFRX1 \block_reg[7][2][9]  ( .D(n1778), .CK(clk), .RN(n3709), .Q(
        \block[7][2][9] ), .QN(n1057) );
  DFFRX1 \block_reg[7][2][8]  ( .D(n1779), .CK(clk), .RN(n3709), .Q(
        \block[7][2][8] ), .QN(n1056) );
  DFFRX1 \block_reg[7][2][7]  ( .D(n1780), .CK(clk), .RN(n3709), .Q(
        \block[7][2][7] ), .QN(n1055) );
  DFFRX1 \block_reg[7][2][6]  ( .D(n1781), .CK(clk), .RN(n3709), .Q(
        \block[7][2][6] ), .QN(n1054) );
  DFFRX1 \block_reg[7][2][5]  ( .D(n1782), .CK(clk), .RN(n3708), .Q(
        \block[7][2][5] ), .QN(n1053) );
  DFFRX1 \block_reg[7][2][4]  ( .D(n1783), .CK(clk), .RN(n3708), .Q(
        \block[7][2][4] ), .QN(n1052) );
  DFFRX1 \block_reg[7][2][3]  ( .D(n1784), .CK(clk), .RN(n3708), .Q(
        \block[7][2][3] ), .QN(n1051) );
  DFFRX1 \block_reg[7][2][2]  ( .D(n1785), .CK(clk), .RN(n3708), .Q(
        \block[7][2][2] ), .QN(n1050) );
  DFFRX1 \block_reg[7][2][1]  ( .D(n1786), .CK(clk), .RN(n3708), .Q(
        \block[7][2][1] ), .QN(n1049) );
  DFFRX1 \block_reg[7][2][0]  ( .D(n1787), .CK(clk), .RN(n3708), .Q(
        \block[7][2][0] ), .QN(n1048) );
  DFFRX1 \block_reg[3][2][31]  ( .D(n2268), .CK(clk), .RN(n3700), .Q(
        \block[3][2][31] ), .QN(n567) );
  DFFRX1 \block_reg[3][2][30]  ( .D(n2269), .CK(clk), .RN(n3700), .Q(
        \block[3][2][30] ), .QN(n566) );
  DFFRX1 \block_reg[3][2][29]  ( .D(n2270), .CK(clk), .RN(n3700), .Q(
        \block[3][2][29] ), .QN(n565) );
  DFFRX1 \block_reg[3][2][28]  ( .D(n2271), .CK(clk), .RN(n3700), .Q(
        \block[3][2][28] ), .QN(n564) );
  DFFRX1 \block_reg[3][2][27]  ( .D(n2272), .CK(clk), .RN(n3700), .Q(
        \block[3][2][27] ), .QN(n563) );
  DFFRX1 \block_reg[3][2][26]  ( .D(n2273), .CK(clk), .RN(n3700), .Q(
        \block[3][2][26] ), .QN(n562) );
  DFFRX1 \block_reg[3][2][25]  ( .D(n2274), .CK(clk), .RN(n3699), .Q(
        \block[3][2][25] ), .QN(n561) );
  DFFRX1 \block_reg[3][2][24]  ( .D(n2275), .CK(clk), .RN(n3699), .Q(
        \block[3][2][24] ), .QN(n560) );
  DFFRX1 \block_reg[3][2][23]  ( .D(n2276), .CK(clk), .RN(n3699), .Q(
        \block[3][2][23] ), .QN(n559) );
  DFFRX1 \block_reg[3][2][22]  ( .D(n2277), .CK(clk), .RN(n3699), .Q(
        \block[3][2][22] ), .QN(n558) );
  DFFRX1 \block_reg[3][2][21]  ( .D(n2278), .CK(clk), .RN(n3699), .Q(
        \block[3][2][21] ), .QN(n557) );
  DFFRX1 \block_reg[3][2][20]  ( .D(n2279), .CK(clk), .RN(n3699), .Q(
        \block[3][2][20] ), .QN(n556) );
  DFFRX1 \block_reg[3][2][19]  ( .D(n2280), .CK(clk), .RN(n3699), .Q(
        \block[3][2][19] ), .QN(n555) );
  DFFRX1 \block_reg[3][2][18]  ( .D(n2281), .CK(clk), .RN(n3699), .Q(
        \block[3][2][18] ), .QN(n554) );
  DFFRX1 \block_reg[3][2][17]  ( .D(n2282), .CK(clk), .RN(n3699), .Q(
        \block[3][2][17] ), .QN(n553) );
  DFFRX1 \block_reg[3][2][16]  ( .D(n2283), .CK(clk), .RN(n3699), .Q(
        \block[3][2][16] ), .QN(n552) );
  DFFRX1 \block_reg[3][2][15]  ( .D(n2284), .CK(clk), .RN(n3699), .Q(
        \block[3][2][15] ), .QN(n551) );
  DFFRX1 \block_reg[3][2][14]  ( .D(n2285), .CK(clk), .RN(n3699), .Q(
        \block[3][2][14] ), .QN(n550) );
  DFFRX1 \block_reg[3][2][13]  ( .D(n2286), .CK(clk), .RN(n3698), .Q(
        \block[3][2][13] ), .QN(n549) );
  DFFRX1 \block_reg[3][2][12]  ( .D(n2287), .CK(clk), .RN(n3698), .Q(
        \block[3][2][12] ), .QN(n548) );
  DFFRX1 \block_reg[3][2][11]  ( .D(n2288), .CK(clk), .RN(n3698), .Q(
        \block[3][2][11] ), .QN(n547) );
  DFFRX1 \block_reg[3][2][10]  ( .D(n2289), .CK(clk), .RN(n3698), .Q(
        \block[3][2][10] ), .QN(n546) );
  DFFRX1 \block_reg[3][2][9]  ( .D(n2290), .CK(clk), .RN(n3698), .Q(
        \block[3][2][9] ), .QN(n545) );
  DFFRX1 \block_reg[3][2][8]  ( .D(n2291), .CK(clk), .RN(n3698), .Q(
        \block[3][2][8] ), .QN(n544) );
  DFFRX1 \block_reg[3][2][7]  ( .D(n2292), .CK(clk), .RN(n3698), .Q(
        \block[3][2][7] ), .QN(n543) );
  DFFRX1 \block_reg[3][2][6]  ( .D(n2293), .CK(clk), .RN(n3698), .Q(
        \block[3][2][6] ), .QN(n542) );
  DFFRX1 \block_reg[3][2][5]  ( .D(n2294), .CK(clk), .RN(n3698), .Q(
        \block[3][2][5] ), .QN(n541) );
  DFFRX1 \block_reg[3][2][4]  ( .D(n2295), .CK(clk), .RN(n3698), .Q(
        \block[3][2][4] ), .QN(n540) );
  DFFRX1 \block_reg[3][2][3]  ( .D(n2296), .CK(clk), .RN(n3698), .Q(
        \block[3][2][3] ), .QN(n539) );
  DFFRX1 \block_reg[3][2][2]  ( .D(n2297), .CK(clk), .RN(n3698), .Q(
        \block[3][2][2] ), .QN(n538) );
  DFFRX1 \block_reg[3][2][1]  ( .D(n2298), .CK(clk), .RN(n3697), .Q(
        \block[3][2][1] ), .QN(n537) );
  DFFRX1 \block_reg[3][2][0]  ( .D(n2299), .CK(clk), .RN(n3697), .Q(
        \block[3][2][0] ), .QN(n536) );
  DFFRX1 \block_reg[7][1][31]  ( .D(n1788), .CK(clk), .RN(n3689), .Q(
        \block[7][1][31] ), .QN(n1047) );
  DFFRX1 \block_reg[7][1][30]  ( .D(n1789), .CK(clk), .RN(n3689), .Q(
        \block[7][1][30] ), .QN(n1046) );
  DFFRX1 \block_reg[7][1][29]  ( .D(n1790), .CK(clk), .RN(n3689), .Q(
        \block[7][1][29] ), .QN(n1045) );
  DFFRX1 \block_reg[7][1][28]  ( .D(n1791), .CK(clk), .RN(n3689), .Q(
        \block[7][1][28] ), .QN(n1044) );
  DFFRX1 \block_reg[7][1][27]  ( .D(n1792), .CK(clk), .RN(n3689), .Q(
        \block[7][1][27] ), .QN(n1043) );
  DFFRX1 \block_reg[7][1][26]  ( .D(n1793), .CK(clk), .RN(n3689), .Q(
        \block[7][1][26] ), .QN(n1042) );
  DFFRX1 \block_reg[7][1][25]  ( .D(n1794), .CK(clk), .RN(n3689), .Q(
        \block[7][1][25] ), .QN(n1041) );
  DFFRX1 \block_reg[7][1][24]  ( .D(n1795), .CK(clk), .RN(n3689), .Q(
        \block[7][1][24] ), .QN(n1040) );
  DFFRX1 \block_reg[7][1][23]  ( .D(n1796), .CK(clk), .RN(n3689), .Q(
        \block[7][1][23] ), .QN(n1039) );
  DFFRX1 \block_reg[7][1][22]  ( .D(n1797), .CK(clk), .RN(n3689), .Q(
        \block[7][1][22] ), .QN(n1038) );
  DFFRX1 \block_reg[7][1][21]  ( .D(n1798), .CK(clk), .RN(n3688), .Q(
        \block[7][1][21] ), .QN(n1037) );
  DFFRX1 \block_reg[7][1][20]  ( .D(n1799), .CK(clk), .RN(n3688), .Q(
        \block[7][1][20] ), .QN(n1036) );
  DFFRX1 \block_reg[7][1][19]  ( .D(n1800), .CK(clk), .RN(n3688), .Q(
        \block[7][1][19] ), .QN(n1035) );
  DFFRX1 \block_reg[7][1][18]  ( .D(n1801), .CK(clk), .RN(n3688), .Q(
        \block[7][1][18] ), .QN(n1034) );
  DFFRX1 \block_reg[7][1][17]  ( .D(n1802), .CK(clk), .RN(n3688), .Q(
        \block[7][1][17] ), .QN(n1033) );
  DFFRX1 \block_reg[7][1][16]  ( .D(n1803), .CK(clk), .RN(n3688), .Q(
        \block[7][1][16] ), .QN(n1032) );
  DFFRX1 \block_reg[7][1][15]  ( .D(n1804), .CK(clk), .RN(n3688), .Q(
        \block[7][1][15] ), .QN(n1031) );
  DFFRX1 \block_reg[7][1][14]  ( .D(n1805), .CK(clk), .RN(n3688), .Q(
        \block[7][1][14] ), .QN(n1030) );
  DFFRX1 \block_reg[7][1][13]  ( .D(n1806), .CK(clk), .RN(n3688), .Q(
        \block[7][1][13] ), .QN(n1029) );
  DFFRX1 \block_reg[7][1][12]  ( .D(n1807), .CK(clk), .RN(n3688), .Q(
        \block[7][1][12] ), .QN(n1028) );
  DFFRX1 \block_reg[7][1][11]  ( .D(n1808), .CK(clk), .RN(n3688), .Q(
        \block[7][1][11] ), .QN(n1027) );
  DFFRX1 \block_reg[7][1][10]  ( .D(n1809), .CK(clk), .RN(n3688), .Q(
        \block[7][1][10] ), .QN(n1026) );
  DFFRX1 \block_reg[7][1][9]  ( .D(n1810), .CK(clk), .RN(n3687), .Q(
        \block[7][1][9] ), .QN(n1025) );
  DFFRX1 \block_reg[7][1][8]  ( .D(n1811), .CK(clk), .RN(n3687), .Q(
        \block[7][1][8] ), .QN(n1024) );
  DFFRX1 \block_reg[7][1][7]  ( .D(n1812), .CK(clk), .RN(n3687), .Q(
        \block[7][1][7] ), .QN(n1023) );
  DFFRX1 \block_reg[7][1][6]  ( .D(n1813), .CK(clk), .RN(n3687), .Q(
        \block[7][1][6] ), .QN(n1022) );
  DFFRX1 \block_reg[7][1][5]  ( .D(n1814), .CK(clk), .RN(n3687), .Q(
        \block[7][1][5] ), .QN(n1021) );
  DFFRX1 \block_reg[7][1][4]  ( .D(n1815), .CK(clk), .RN(n3687), .Q(
        \block[7][1][4] ), .QN(n1020) );
  DFFRX1 \block_reg[7][1][3]  ( .D(n1816), .CK(clk), .RN(n3687), .Q(
        \block[7][1][3] ), .QN(n1019) );
  DFFRX1 \block_reg[7][1][2]  ( .D(n1817), .CK(clk), .RN(n3687), .Q(
        \block[7][1][2] ), .QN(n1018) );
  DFFRX1 \block_reg[7][1][1]  ( .D(n1818), .CK(clk), .RN(n3687), .Q(
        \block[7][1][1] ), .QN(n1017) );
  DFFRX1 \block_reg[7][1][0]  ( .D(n1819), .CK(clk), .RN(n3687), .Q(
        \block[7][1][0] ), .QN(n1016) );
  DFFRX1 \block_reg[3][1][31]  ( .D(n2300), .CK(clk), .RN(n3679), .Q(
        \block[3][1][31] ), .QN(n535) );
  DFFRX1 \block_reg[3][1][30]  ( .D(n2301), .CK(clk), .RN(n3679), .Q(
        \block[3][1][30] ), .QN(n534) );
  DFFRX1 \block_reg[3][1][29]  ( .D(n2302), .CK(clk), .RN(n3678), .Q(
        \block[3][1][29] ), .QN(n533) );
  DFFRX1 \block_reg[3][1][28]  ( .D(n2303), .CK(clk), .RN(n3678), .Q(
        \block[3][1][28] ), .QN(n532) );
  DFFRX1 \block_reg[3][1][27]  ( .D(n2304), .CK(clk), .RN(n3678), .Q(
        \block[3][1][27] ), .QN(n531) );
  DFFRX1 \block_reg[3][1][26]  ( .D(n2305), .CK(clk), .RN(n3678), .Q(
        \block[3][1][26] ), .QN(n530) );
  DFFRX1 \block_reg[3][1][25]  ( .D(n2306), .CK(clk), .RN(n3678), .Q(
        \block[3][1][25] ), .QN(n529) );
  DFFRX1 \block_reg[3][1][24]  ( .D(n2307), .CK(clk), .RN(n3678), .Q(
        \block[3][1][24] ), .QN(n528) );
  DFFRX1 \block_reg[3][1][23]  ( .D(n2308), .CK(clk), .RN(n3678), .Q(
        \block[3][1][23] ), .QN(n527) );
  DFFRX1 \block_reg[3][1][22]  ( .D(n2309), .CK(clk), .RN(n3678), .Q(
        \block[3][1][22] ), .QN(n526) );
  DFFRX1 \block_reg[3][1][21]  ( .D(n2310), .CK(clk), .RN(n3678), .Q(
        \block[3][1][21] ), .QN(n525) );
  DFFRX1 \block_reg[3][1][20]  ( .D(n2311), .CK(clk), .RN(n3678), .Q(
        \block[3][1][20] ), .QN(n524) );
  DFFRX1 \block_reg[3][1][19]  ( .D(n2312), .CK(clk), .RN(n3678), .Q(
        \block[3][1][19] ), .QN(n523) );
  DFFRX1 \block_reg[3][1][18]  ( .D(n2313), .CK(clk), .RN(n3678), .Q(
        \block[3][1][18] ), .QN(n522) );
  DFFRX1 \block_reg[3][1][17]  ( .D(n2314), .CK(clk), .RN(n3677), .Q(
        \block[3][1][17] ), .QN(n521) );
  DFFRX1 \block_reg[3][1][16]  ( .D(n2315), .CK(clk), .RN(n3677), .Q(
        \block[3][1][16] ), .QN(n520) );
  DFFRX1 \block_reg[3][1][15]  ( .D(n2316), .CK(clk), .RN(n3677), .Q(
        \block[3][1][15] ), .QN(n519) );
  DFFRX1 \block_reg[3][1][14]  ( .D(n2317), .CK(clk), .RN(n3677), .Q(
        \block[3][1][14] ), .QN(n518) );
  DFFRX1 \block_reg[3][1][13]  ( .D(n2318), .CK(clk), .RN(n3677), .Q(
        \block[3][1][13] ), .QN(n517) );
  DFFRX1 \block_reg[3][1][12]  ( .D(n2319), .CK(clk), .RN(n3677), .Q(
        \block[3][1][12] ), .QN(n516) );
  DFFRX1 \block_reg[3][1][11]  ( .D(n2320), .CK(clk), .RN(n3677), .Q(
        \block[3][1][11] ), .QN(n515) );
  DFFRX1 \block_reg[3][1][10]  ( .D(n2321), .CK(clk), .RN(n3677), .Q(
        \block[3][1][10] ), .QN(n514) );
  DFFRX1 \block_reg[3][1][9]  ( .D(n2322), .CK(clk), .RN(n3677), .Q(
        \block[3][1][9] ), .QN(n513) );
  DFFRX1 \block_reg[3][1][8]  ( .D(n2323), .CK(clk), .RN(n3677), .Q(
        \block[3][1][8] ), .QN(n512) );
  DFFRX1 \block_reg[3][1][7]  ( .D(n2324), .CK(clk), .RN(n3677), .Q(
        \block[3][1][7] ), .QN(n511) );
  DFFRX1 \block_reg[3][1][6]  ( .D(n2325), .CK(clk), .RN(n3677), .Q(
        \block[3][1][6] ), .QN(n510) );
  DFFRX1 \block_reg[3][1][5]  ( .D(n2326), .CK(clk), .RN(n3676), .Q(
        \block[3][1][5] ), .QN(n509) );
  DFFRX1 \block_reg[3][1][4]  ( .D(n2327), .CK(clk), .RN(n3676), .Q(
        \block[3][1][4] ), .QN(n508) );
  DFFRX1 \block_reg[3][1][3]  ( .D(n2328), .CK(clk), .RN(n3676), .Q(
        \block[3][1][3] ), .QN(n507) );
  DFFRX1 \block_reg[3][1][2]  ( .D(n2329), .CK(clk), .RN(n3676), .Q(
        \block[3][1][2] ), .QN(n506) );
  DFFRX1 \block_reg[3][1][1]  ( .D(n2330), .CK(clk), .RN(n3676), .Q(
        \block[3][1][1] ), .QN(n505) );
  DFFRX1 \block_reg[3][1][0]  ( .D(n2331), .CK(clk), .RN(n3676), .Q(
        \block[3][1][0] ), .QN(n504) );
  DFFRX1 \block_reg[2][0][31]  ( .D(n2460), .CK(clk), .RN(n3759), .Q(
        \block[2][0][31] ), .QN(n1670) );
  DFFRX1 \block_reg[2][0][30]  ( .D(n2461), .CK(clk), .RN(n3759), .Q(
        \block[2][0][30] ), .QN(n1669) );
  DFFRX1 \block_reg[2][0][29]  ( .D(n2462), .CK(clk), .RN(n3758), .Q(
        \block[2][0][29] ), .QN(n1668) );
  DFFRX1 \block_reg[2][0][28]  ( .D(n2463), .CK(clk), .RN(n3758), .Q(
        \block[2][0][28] ), .QN(n1667) );
  DFFRX1 \block_reg[2][0][27]  ( .D(n2464), .CK(clk), .RN(n3758), .Q(
        \block[2][0][27] ), .QN(n1666) );
  DFFRX1 \block_reg[2][0][26]  ( .D(n2465), .CK(clk), .RN(n3758), .Q(
        \block[2][0][26] ), .QN(n1665) );
  DFFRX1 \block_reg[2][0][25]  ( .D(n2466), .CK(clk), .RN(n3758), .Q(
        \block[2][0][25] ), .QN(n1664) );
  DFFRX1 \block_reg[2][0][24]  ( .D(n2467), .CK(clk), .RN(n3758), .Q(
        \block[2][0][24] ), .QN(n1663) );
  DFFRX1 \block_reg[2][0][23]  ( .D(n2468), .CK(clk), .RN(n3758), .Q(
        \block[2][0][23] ), .QN(n1662) );
  DFFRX1 \block_reg[2][0][22]  ( .D(n2469), .CK(clk), .RN(n3758), .Q(
        \block[2][0][22] ), .QN(n1661) );
  DFFRX1 \block_reg[2][0][21]  ( .D(n2470), .CK(clk), .RN(n3758), .Q(
        \block[2][0][21] ), .QN(n1660) );
  DFFRX1 \block_reg[2][0][20]  ( .D(n2471), .CK(clk), .RN(n3758), .Q(
        \block[2][0][20] ), .QN(n1659) );
  DFFRX1 \block_reg[2][0][19]  ( .D(n2472), .CK(clk), .RN(n3758), .Q(
        \block[2][0][19] ), .QN(n1658) );
  DFFRX1 \block_reg[2][0][18]  ( .D(n2473), .CK(clk), .RN(n3758), .Q(
        \block[2][0][18] ), .QN(n1657) );
  DFFRX1 \block_reg[2][0][17]  ( .D(n2474), .CK(clk), .RN(n3757), .Q(
        \block[2][0][17] ), .QN(n1656) );
  DFFRX1 \block_reg[2][0][16]  ( .D(n2475), .CK(clk), .RN(n3757), .Q(
        \block[2][0][16] ), .QN(n1655) );
  DFFRX1 \block_reg[2][0][15]  ( .D(n2476), .CK(clk), .RN(n3757), .Q(
        \block[2][0][15] ), .QN(n1654) );
  DFFRX1 \block_reg[2][0][14]  ( .D(n2477), .CK(clk), .RN(n3757), .Q(
        \block[2][0][14] ), .QN(n1653) );
  DFFRX1 \block_reg[2][0][13]  ( .D(n2478), .CK(clk), .RN(n3757), .Q(
        \block[2][0][13] ), .QN(n1652) );
  DFFRX1 \block_reg[2][0][12]  ( .D(n2479), .CK(clk), .RN(n3757), .Q(
        \block[2][0][12] ), .QN(n1651) );
  DFFRX1 \block_reg[2][0][11]  ( .D(n2480), .CK(clk), .RN(n3757), .Q(
        \block[2][0][11] ), .QN(n1650) );
  DFFRX1 \block_reg[2][0][10]  ( .D(n2481), .CK(clk), .RN(n3757), .Q(
        \block[2][0][10] ), .QN(n1649) );
  DFFRX1 \block_reg[2][0][9]  ( .D(n2482), .CK(clk), .RN(n3757), .Q(
        \block[2][0][9] ), .QN(n1648) );
  DFFRX1 \block_reg[2][0][8]  ( .D(n2483), .CK(clk), .RN(n3757), .Q(
        \block[2][0][8] ), .QN(n1647) );
  DFFRX1 \block_reg[2][0][7]  ( .D(n2484), .CK(clk), .RN(n3757), .Q(
        \block[2][0][7] ), .QN(n1646) );
  DFFRX1 \block_reg[2][0][6]  ( .D(n2485), .CK(clk), .RN(n3757), .Q(
        \block[2][0][6] ), .QN(n1645) );
  DFFRX1 \block_reg[2][0][5]  ( .D(n2486), .CK(clk), .RN(n3756), .Q(
        \block[2][0][5] ), .QN(n1644) );
  DFFRX1 \block_reg[2][0][4]  ( .D(n2487), .CK(clk), .RN(n3756), .Q(
        \block[2][0][4] ), .QN(n1643) );
  DFFRX1 \block_reg[2][0][3]  ( .D(n2488), .CK(clk), .RN(n3756), .Q(
        \block[2][0][3] ), .QN(n1642) );
  DFFRX1 \block_reg[2][0][2]  ( .D(n2489), .CK(clk), .RN(n3756), .Q(
        \block[2][0][2] ), .QN(n1641) );
  DFFRX1 \block_reg[2][0][1]  ( .D(n2490), .CK(clk), .RN(n3756), .Q(
        \block[2][0][1] ), .QN(n1640) );
  DFFRX1 \block_reg[2][0][0]  ( .D(n2491), .CK(clk), .RN(n3756), .Q(
        \block[2][0][0] ), .QN(n1639) );
  DFFRX1 \block_reg[6][0][31]  ( .D(n1948), .CK(clk), .RN(n3748), .Q(
        \block[6][0][31] ), .QN(n887) );
  DFFRX1 \block_reg[6][0][30]  ( .D(n1949), .CK(clk), .RN(n3748), .Q(
        \block[6][0][30] ), .QN(n886) );
  DFFRX1 \block_reg[6][0][29]  ( .D(n1950), .CK(clk), .RN(n3748), .Q(
        \block[6][0][29] ), .QN(n885) );
  DFFRX1 \block_reg[6][0][28]  ( .D(n1951), .CK(clk), .RN(n3748), .Q(
        \block[6][0][28] ), .QN(n884) );
  DFFRX1 \block_reg[6][0][27]  ( .D(n1952), .CK(clk), .RN(n3748), .Q(
        \block[6][0][27] ), .QN(n883) );
  DFFRX1 \block_reg[6][0][26]  ( .D(n1953), .CK(clk), .RN(n3748), .Q(
        \block[6][0][26] ), .QN(n882) );
  DFFRX1 \block_reg[6][0][25]  ( .D(n1954), .CK(clk), .RN(n3747), .Q(
        \block[6][0][25] ), .QN(n881) );
  DFFRX1 \block_reg[6][0][24]  ( .D(n1955), .CK(clk), .RN(n3747), .Q(
        \block[6][0][24] ), .QN(n880) );
  DFFRX1 \block_reg[6][0][23]  ( .D(n1956), .CK(clk), .RN(n3747), .Q(
        \block[6][0][23] ), .QN(n879) );
  DFFRX1 \block_reg[6][0][22]  ( .D(n1957), .CK(clk), .RN(n3747), .Q(
        \block[6][0][22] ), .QN(n878) );
  DFFRX1 \block_reg[6][0][21]  ( .D(n1958), .CK(clk), .RN(n3747), .Q(
        \block[6][0][21] ), .QN(n877) );
  DFFRX1 \block_reg[6][0][20]  ( .D(n1959), .CK(clk), .RN(n3747), .Q(
        \block[6][0][20] ), .QN(n876) );
  DFFRX1 \block_reg[6][0][19]  ( .D(n1960), .CK(clk), .RN(n3747), .Q(
        \block[6][0][19] ), .QN(n875) );
  DFFRX1 \block_reg[6][0][18]  ( .D(n1961), .CK(clk), .RN(n3747), .Q(
        \block[6][0][18] ), .QN(n874) );
  DFFRX1 \block_reg[6][0][17]  ( .D(n1962), .CK(clk), .RN(n3747), .Q(
        \block[6][0][17] ), .QN(n873) );
  DFFRX1 \block_reg[6][0][16]  ( .D(n1963), .CK(clk), .RN(n3747), .Q(
        \block[6][0][16] ), .QN(n872) );
  DFFRX1 \block_reg[6][0][15]  ( .D(n1964), .CK(clk), .RN(n3747), .Q(
        \block[6][0][15] ), .QN(n871) );
  DFFRX1 \block_reg[6][0][14]  ( .D(n1965), .CK(clk), .RN(n3747), .Q(
        \block[6][0][14] ), .QN(n870) );
  DFFRX1 \block_reg[6][0][13]  ( .D(n1966), .CK(clk), .RN(n3746), .Q(
        \block[6][0][13] ), .QN(n869) );
  DFFRX1 \block_reg[6][0][12]  ( .D(n1967), .CK(clk), .RN(n3746), .Q(
        \block[6][0][12] ), .QN(n868) );
  DFFRX1 \block_reg[6][0][11]  ( .D(n1968), .CK(clk), .RN(n3746), .Q(
        \block[6][0][11] ), .QN(n867) );
  DFFRX1 \block_reg[6][0][10]  ( .D(n1969), .CK(clk), .RN(n3746), .Q(
        \block[6][0][10] ), .QN(n866) );
  DFFRX1 \block_reg[6][0][9]  ( .D(n1970), .CK(clk), .RN(n3746), .Q(
        \block[6][0][9] ), .QN(n865) );
  DFFRX1 \block_reg[6][0][8]  ( .D(n1971), .CK(clk), .RN(n3746), .Q(
        \block[6][0][8] ), .QN(n864) );
  DFFRX1 \block_reg[6][0][7]  ( .D(n1972), .CK(clk), .RN(n3746), .Q(
        \block[6][0][7] ), .QN(n863) );
  DFFRX1 \block_reg[6][0][6]  ( .D(n1973), .CK(clk), .RN(n3746), .Q(
        \block[6][0][6] ), .QN(n862) );
  DFFRX1 \block_reg[6][0][5]  ( .D(n1974), .CK(clk), .RN(n3746), .Q(
        \block[6][0][5] ), .QN(n861) );
  DFFRX1 \block_reg[6][0][4]  ( .D(n1975), .CK(clk), .RN(n3746), .Q(
        \block[6][0][4] ), .QN(n860) );
  DFFRX1 \block_reg[6][0][3]  ( .D(n1976), .CK(clk), .RN(n3746), .Q(
        \block[6][0][3] ), .QN(n859) );
  DFFRX1 \block_reg[6][0][2]  ( .D(n1977), .CK(clk), .RN(n3746), .Q(
        \block[6][0][2] ), .QN(n858) );
  DFFRX1 \block_reg[6][0][1]  ( .D(n1978), .CK(clk), .RN(n3745), .Q(
        \block[6][0][1] ), .QN(n857) );
  DFFRX1 \block_reg[6][0][0]  ( .D(n1979), .CK(clk), .RN(n3745), .Q(
        \block[6][0][0] ), .QN(n856) );
  DFFRX1 \block_reg[6][3][31]  ( .D(n1852), .CK(clk), .RN(n3729), .Q(
        \block[6][3][31] ), .QN(n983) );
  DFFRX1 \block_reg[6][3][30]  ( .D(n1853), .CK(clk), .RN(n3729), .Q(
        \block[6][3][30] ), .QN(n982) );
  DFFRX1 \block_reg[6][3][29]  ( .D(n1854), .CK(clk), .RN(n3729), .Q(
        \block[6][3][29] ), .QN(n981) );
  DFFRX1 \block_reg[6][3][28]  ( .D(n1855), .CK(clk), .RN(n3729), .Q(
        \block[6][3][28] ), .QN(n980) );
  DFFRX1 \block_reg[6][3][27]  ( .D(n1856), .CK(clk), .RN(n3729), .Q(
        \block[6][3][27] ), .QN(n979) );
  DFFRX1 \block_reg[6][3][26]  ( .D(n1857), .CK(clk), .RN(n3729), .Q(
        \block[6][3][26] ), .QN(n978) );
  DFFRX1 \block_reg[6][3][25]  ( .D(n1858), .CK(clk), .RN(n3729), .Q(
        \block[6][3][25] ), .QN(n977) );
  DFFRX1 \block_reg[6][3][24]  ( .D(n1859), .CK(clk), .RN(n3729), .Q(
        \block[6][3][24] ), .QN(n976) );
  DFFRX1 \block_reg[6][3][23]  ( .D(n1860), .CK(clk), .RN(n3729), .Q(
        \block[6][3][23] ), .QN(n975) );
  DFFRX1 \block_reg[6][3][22]  ( .D(n1861), .CK(clk), .RN(n3729), .Q(
        \block[6][3][22] ), .QN(n974) );
  DFFRX1 \block_reg[6][3][21]  ( .D(n1862), .CK(clk), .RN(n3728), .Q(
        \block[6][3][21] ), .QN(n973) );
  DFFRX1 \block_reg[6][3][20]  ( .D(n1863), .CK(clk), .RN(n3728), .Q(
        \block[6][3][20] ), .QN(n972) );
  DFFRX1 \block_reg[6][3][19]  ( .D(n1864), .CK(clk), .RN(n3728), .Q(
        \block[6][3][19] ), .QN(n971) );
  DFFRX1 \block_reg[6][3][18]  ( .D(n1865), .CK(clk), .RN(n3728), .Q(
        \block[6][3][18] ), .QN(n970) );
  DFFRX1 \block_reg[6][3][17]  ( .D(n1866), .CK(clk), .RN(n3728), .Q(
        \block[6][3][17] ), .QN(n969) );
  DFFRX1 \block_reg[6][3][16]  ( .D(n1867), .CK(clk), .RN(n3728), .Q(
        \block[6][3][16] ), .QN(n968) );
  DFFRX1 \block_reg[6][3][15]  ( .D(n1868), .CK(clk), .RN(n3728), .Q(
        \block[6][3][15] ), .QN(n967) );
  DFFRX1 \block_reg[6][3][14]  ( .D(n1869), .CK(clk), .RN(n3728), .Q(
        \block[6][3][14] ), .QN(n966) );
  DFFRX1 \block_reg[6][3][13]  ( .D(n1870), .CK(clk), .RN(n3728), .Q(
        \block[6][3][13] ), .QN(n965) );
  DFFRX1 \block_reg[6][3][12]  ( .D(n1871), .CK(clk), .RN(n3728), .Q(
        \block[6][3][12] ), .QN(n964) );
  DFFRX1 \block_reg[6][3][11]  ( .D(n1872), .CK(clk), .RN(n3728), .Q(
        \block[6][3][11] ), .QN(n963) );
  DFFRX1 \block_reg[6][3][10]  ( .D(n1873), .CK(clk), .RN(n3728), .Q(
        \block[6][3][10] ), .QN(n962) );
  DFFRX1 \block_reg[6][3][9]  ( .D(n1874), .CK(clk), .RN(n3727), .Q(
        \block[6][3][9] ), .QN(n961) );
  DFFRX1 \block_reg[6][3][8]  ( .D(n1875), .CK(clk), .RN(n3727), .Q(
        \block[6][3][8] ), .QN(n960) );
  DFFRX1 \block_reg[6][3][7]  ( .D(n1876), .CK(clk), .RN(n3727), .Q(
        \block[6][3][7] ), .QN(n959) );
  DFFRX1 \block_reg[6][3][6]  ( .D(n1877), .CK(clk), .RN(n3727), .Q(
        \block[6][3][6] ), .QN(n958) );
  DFFRX1 \block_reg[6][3][5]  ( .D(n1878), .CK(clk), .RN(n3727), .Q(
        \block[6][3][5] ), .QN(n957) );
  DFFRX1 \block_reg[6][3][4]  ( .D(n1879), .CK(clk), .RN(n3727), .Q(
        \block[6][3][4] ), .QN(n956) );
  DFFRX1 \block_reg[6][3][3]  ( .D(n1880), .CK(clk), .RN(n3727), .Q(
        \block[6][3][3] ), .QN(n955) );
  DFFRX1 \block_reg[6][3][2]  ( .D(n1881), .CK(clk), .RN(n3727), .Q(
        \block[6][3][2] ), .QN(n954) );
  DFFRX1 \block_reg[6][3][1]  ( .D(n1882), .CK(clk), .RN(n3727), .Q(
        \block[6][3][1] ), .QN(n953) );
  DFFRX1 \block_reg[6][3][0]  ( .D(n1883), .CK(clk), .RN(n3727), .Q(
        \block[6][3][0] ), .QN(n952) );
  DFFRX1 \block_reg[2][3][31]  ( .D(n2364), .CK(clk), .RN(n3719), .Q(
        \block[2][3][31] ), .QN(n471) );
  DFFRX1 \block_reg[2][3][30]  ( .D(n2365), .CK(clk), .RN(n3719), .Q(
        \block[2][3][30] ), .QN(n470) );
  DFFRX1 \block_reg[2][3][29]  ( .D(n2366), .CK(clk), .RN(n3718), .Q(
        \block[2][3][29] ), .QN(n469) );
  DFFRX1 \block_reg[2][3][28]  ( .D(n2367), .CK(clk), .RN(n3718), .Q(
        \block[2][3][28] ), .QN(n468) );
  DFFRX1 \block_reg[2][3][27]  ( .D(n2368), .CK(clk), .RN(n3718), .Q(
        \block[2][3][27] ), .QN(n467) );
  DFFRX1 \block_reg[2][3][26]  ( .D(n2369), .CK(clk), .RN(n3718), .Q(
        \block[2][3][26] ), .QN(n466) );
  DFFRX1 \block_reg[2][3][25]  ( .D(n2370), .CK(clk), .RN(n3718), .Q(
        \block[2][3][25] ), .QN(n465) );
  DFFRX1 \block_reg[2][3][24]  ( .D(n2371), .CK(clk), .RN(n3718), .Q(
        \block[2][3][24] ), .QN(n464) );
  DFFRX1 \block_reg[2][3][23]  ( .D(n2372), .CK(clk), .RN(n3718), .Q(
        \block[2][3][23] ), .QN(n463) );
  DFFRX1 \block_reg[2][3][22]  ( .D(n2373), .CK(clk), .RN(n3718), .Q(
        \block[2][3][22] ), .QN(n462) );
  DFFRX1 \block_reg[2][3][21]  ( .D(n2374), .CK(clk), .RN(n3718), .Q(
        \block[2][3][21] ), .QN(n461) );
  DFFRX1 \block_reg[2][3][20]  ( .D(n2375), .CK(clk), .RN(n3718), .Q(
        \block[2][3][20] ), .QN(n460) );
  DFFRX1 \block_reg[2][3][19]  ( .D(n2376), .CK(clk), .RN(n3718), .Q(
        \block[2][3][19] ), .QN(n459) );
  DFFRX1 \block_reg[2][3][18]  ( .D(n2377), .CK(clk), .RN(n3718), .Q(
        \block[2][3][18] ), .QN(n458) );
  DFFRX1 \block_reg[2][3][17]  ( .D(n2378), .CK(clk), .RN(n3717), .Q(
        \block[2][3][17] ), .QN(n457) );
  DFFRX1 \block_reg[2][3][16]  ( .D(n2379), .CK(clk), .RN(n3717), .Q(
        \block[2][3][16] ), .QN(n456) );
  DFFRX1 \block_reg[2][3][15]  ( .D(n2380), .CK(clk), .RN(n3717), .Q(
        \block[2][3][15] ), .QN(n455) );
  DFFRX1 \block_reg[2][3][14]  ( .D(n2381), .CK(clk), .RN(n3717), .Q(
        \block[2][3][14] ), .QN(n454) );
  DFFRX1 \block_reg[2][3][13]  ( .D(n2382), .CK(clk), .RN(n3717), .Q(
        \block[2][3][13] ), .QN(n453) );
  DFFRX1 \block_reg[2][3][12]  ( .D(n2383), .CK(clk), .RN(n3717), .Q(
        \block[2][3][12] ), .QN(n452) );
  DFFRX1 \block_reg[2][3][11]  ( .D(n2384), .CK(clk), .RN(n3717), .Q(
        \block[2][3][11] ), .QN(n451) );
  DFFRX1 \block_reg[2][3][10]  ( .D(n2385), .CK(clk), .RN(n3717), .Q(
        \block[2][3][10] ), .QN(n450) );
  DFFRX1 \block_reg[2][3][9]  ( .D(n2386), .CK(clk), .RN(n3717), .Q(
        \block[2][3][9] ), .QN(n449) );
  DFFRX1 \block_reg[2][3][8]  ( .D(n2387), .CK(clk), .RN(n3717), .Q(
        \block[2][3][8] ), .QN(n448) );
  DFFRX1 \block_reg[2][3][7]  ( .D(n2388), .CK(clk), .RN(n3717), .Q(
        \block[2][3][7] ), .QN(n447) );
  DFFRX1 \block_reg[2][3][6]  ( .D(n2389), .CK(clk), .RN(n3717), .Q(
        \block[2][3][6] ), .QN(n446) );
  DFFRX1 \block_reg[2][3][5]  ( .D(n2390), .CK(clk), .RN(n3716), .Q(
        \block[2][3][5] ), .QN(n445) );
  DFFRX1 \block_reg[2][3][4]  ( .D(n2391), .CK(clk), .RN(n3716), .Q(
        \block[2][3][4] ), .QN(n444) );
  DFFRX1 \block_reg[2][3][3]  ( .D(n2392), .CK(clk), .RN(n3716), .Q(
        \block[2][3][3] ), .QN(n443) );
  DFFRX1 \block_reg[2][3][2]  ( .D(n2393), .CK(clk), .RN(n3716), .Q(
        \block[2][3][2] ), .QN(n442) );
  DFFRX1 \block_reg[2][3][1]  ( .D(n2394), .CK(clk), .RN(n3716), .Q(
        \block[2][3][1] ), .QN(n441) );
  DFFRX1 \block_reg[2][3][0]  ( .D(n2395), .CK(clk), .RN(n3716), .Q(
        \block[2][3][0] ), .QN(n440) );
  DFFRX1 \block_reg[6][2][31]  ( .D(n1884), .CK(clk), .RN(n3708), .Q(
        \block[6][2][31] ), .QN(n951) );
  DFFRX1 \block_reg[6][2][30]  ( .D(n1885), .CK(clk), .RN(n3708), .Q(
        \block[6][2][30] ), .QN(n950) );
  DFFRX1 \block_reg[6][2][29]  ( .D(n1886), .CK(clk), .RN(n3708), .Q(
        \block[6][2][29] ), .QN(n949) );
  DFFRX1 \block_reg[6][2][28]  ( .D(n1887), .CK(clk), .RN(n3708), .Q(
        \block[6][2][28] ), .QN(n948) );
  DFFRX1 \block_reg[6][2][27]  ( .D(n1888), .CK(clk), .RN(n3708), .Q(
        \block[6][2][27] ), .QN(n947) );
  DFFRX1 \block_reg[6][2][26]  ( .D(n1889), .CK(clk), .RN(n3708), .Q(
        \block[6][2][26] ), .QN(n946) );
  DFFRX1 \block_reg[6][2][25]  ( .D(n1890), .CK(clk), .RN(n3707), .Q(
        \block[6][2][25] ), .QN(n945) );
  DFFRX1 \block_reg[6][2][24]  ( .D(n1891), .CK(clk), .RN(n3707), .Q(
        \block[6][2][24] ), .QN(n944) );
  DFFRX1 \block_reg[6][2][23]  ( .D(n1892), .CK(clk), .RN(n3707), .Q(
        \block[6][2][23] ), .QN(n943) );
  DFFRX1 \block_reg[6][2][22]  ( .D(n1893), .CK(clk), .RN(n3707), .Q(
        \block[6][2][22] ), .QN(n942) );
  DFFRX1 \block_reg[6][2][21]  ( .D(n1894), .CK(clk), .RN(n3707), .Q(
        \block[6][2][21] ), .QN(n941) );
  DFFRX1 \block_reg[6][2][20]  ( .D(n1895), .CK(clk), .RN(n3707), .Q(
        \block[6][2][20] ), .QN(n940) );
  DFFRX1 \block_reg[6][2][19]  ( .D(n1896), .CK(clk), .RN(n3707), .Q(
        \block[6][2][19] ), .QN(n939) );
  DFFRX1 \block_reg[6][2][18]  ( .D(n1897), .CK(clk), .RN(n3707), .Q(
        \block[6][2][18] ), .QN(n938) );
  DFFRX1 \block_reg[6][2][17]  ( .D(n1898), .CK(clk), .RN(n3707), .Q(
        \block[6][2][17] ), .QN(n937) );
  DFFRX1 \block_reg[6][2][16]  ( .D(n1899), .CK(clk), .RN(n3707), .Q(
        \block[6][2][16] ), .QN(n936) );
  DFFRX1 \block_reg[6][2][15]  ( .D(n1900), .CK(clk), .RN(n3707), .Q(
        \block[6][2][15] ), .QN(n935) );
  DFFRX1 \block_reg[6][2][14]  ( .D(n1901), .CK(clk), .RN(n3707), .Q(
        \block[6][2][14] ), .QN(n934) );
  DFFRX1 \block_reg[6][2][13]  ( .D(n1902), .CK(clk), .RN(n3706), .Q(
        \block[6][2][13] ), .QN(n933) );
  DFFRX1 \block_reg[6][2][12]  ( .D(n1903), .CK(clk), .RN(n3706), .Q(
        \block[6][2][12] ), .QN(n932) );
  DFFRX1 \block_reg[6][2][11]  ( .D(n1904), .CK(clk), .RN(n3706), .Q(
        \block[6][2][11] ), .QN(n931) );
  DFFRX1 \block_reg[6][2][10]  ( .D(n1905), .CK(clk), .RN(n3706), .Q(
        \block[6][2][10] ), .QN(n930) );
  DFFRX1 \block_reg[6][2][9]  ( .D(n1906), .CK(clk), .RN(n3706), .Q(
        \block[6][2][9] ), .QN(n929) );
  DFFRX1 \block_reg[6][2][8]  ( .D(n1907), .CK(clk), .RN(n3706), .Q(
        \block[6][2][8] ), .QN(n928) );
  DFFRX1 \block_reg[6][2][7]  ( .D(n1908), .CK(clk), .RN(n3706), .Q(
        \block[6][2][7] ), .QN(n927) );
  DFFRX1 \block_reg[6][2][6]  ( .D(n1909), .CK(clk), .RN(n3706), .Q(
        \block[6][2][6] ), .QN(n926) );
  DFFRX1 \block_reg[6][2][5]  ( .D(n1910), .CK(clk), .RN(n3706), .Q(
        \block[6][2][5] ), .QN(n925) );
  DFFRX1 \block_reg[6][2][4]  ( .D(n1911), .CK(clk), .RN(n3706), .Q(
        \block[6][2][4] ), .QN(n924) );
  DFFRX1 \block_reg[6][2][3]  ( .D(n1912), .CK(clk), .RN(n3706), .Q(
        \block[6][2][3] ), .QN(n923) );
  DFFRX1 \block_reg[6][2][2]  ( .D(n1913), .CK(clk), .RN(n3706), .Q(
        \block[6][2][2] ), .QN(n922) );
  DFFRX1 \block_reg[6][2][1]  ( .D(n1914), .CK(clk), .RN(n3705), .Q(
        \block[6][2][1] ), .QN(n921) );
  DFFRX1 \block_reg[6][2][0]  ( .D(n1915), .CK(clk), .RN(n3705), .Q(
        \block[6][2][0] ), .QN(n920) );
  DFFRX1 \block_reg[2][2][31]  ( .D(n2396), .CK(clk), .RN(n3697), .Q(
        \block[2][2][31] ), .QN(n439) );
  DFFRX1 \block_reg[2][2][30]  ( .D(n2397), .CK(clk), .RN(n3697), .Q(
        \block[2][2][30] ), .QN(n438) );
  DFFRX1 \block_reg[2][2][29]  ( .D(n2398), .CK(clk), .RN(n3697), .Q(
        \block[2][2][29] ), .QN(n437) );
  DFFRX1 \block_reg[2][2][28]  ( .D(n2399), .CK(clk), .RN(n3697), .Q(
        \block[2][2][28] ), .QN(n436) );
  DFFRX1 \block_reg[2][2][27]  ( .D(n2400), .CK(clk), .RN(n3697), .Q(
        \block[2][2][27] ), .QN(n435) );
  DFFRX1 \block_reg[2][2][26]  ( .D(n2401), .CK(clk), .RN(n3697), .Q(
        \block[2][2][26] ), .QN(n434) );
  DFFRX1 \block_reg[2][2][25]  ( .D(n2402), .CK(clk), .RN(n3697), .Q(
        \block[2][2][25] ), .QN(n433) );
  DFFRX1 \block_reg[2][2][24]  ( .D(n2403), .CK(clk), .RN(n3697), .Q(
        \block[2][2][24] ), .QN(n432) );
  DFFRX1 \block_reg[2][2][23]  ( .D(n2404), .CK(clk), .RN(n3697), .Q(
        \block[2][2][23] ), .QN(n431) );
  DFFRX1 \block_reg[2][2][22]  ( .D(n2405), .CK(clk), .RN(n3697), .Q(
        \block[2][2][22] ), .QN(n430) );
  DFFRX1 \block_reg[2][2][21]  ( .D(n2406), .CK(clk), .RN(n3696), .Q(
        \block[2][2][21] ), .QN(n429) );
  DFFRX1 \block_reg[2][2][20]  ( .D(n2407), .CK(clk), .RN(n3696), .Q(
        \block[2][2][20] ), .QN(n428) );
  DFFRX1 \block_reg[2][2][19]  ( .D(n2408), .CK(clk), .RN(n3696), .Q(
        \block[2][2][19] ), .QN(n427) );
  DFFRX1 \block_reg[2][2][18]  ( .D(n2409), .CK(clk), .RN(n3696), .Q(
        \block[2][2][18] ), .QN(n426) );
  DFFRX1 \block_reg[2][2][17]  ( .D(n2410), .CK(clk), .RN(n3696), .Q(
        \block[2][2][17] ), .QN(n425) );
  DFFRX1 \block_reg[2][2][16]  ( .D(n2411), .CK(clk), .RN(n3696), .Q(
        \block[2][2][16] ), .QN(n424) );
  DFFRX1 \block_reg[2][2][15]  ( .D(n2412), .CK(clk), .RN(n3696), .Q(
        \block[2][2][15] ), .QN(n423) );
  DFFRX1 \block_reg[2][2][14]  ( .D(n2413), .CK(clk), .RN(n3696), .Q(
        \block[2][2][14] ), .QN(n422) );
  DFFRX1 \block_reg[2][2][13]  ( .D(n2414), .CK(clk), .RN(n3696), .Q(
        \block[2][2][13] ), .QN(n421) );
  DFFRX1 \block_reg[2][2][12]  ( .D(n2415), .CK(clk), .RN(n3696), .Q(
        \block[2][2][12] ), .QN(n420) );
  DFFRX1 \block_reg[2][2][11]  ( .D(n2416), .CK(clk), .RN(n3696), .Q(
        \block[2][2][11] ), .QN(n419) );
  DFFRX1 \block_reg[2][2][10]  ( .D(n2417), .CK(clk), .RN(n3696), .Q(
        \block[2][2][10] ), .QN(n418) );
  DFFRX1 \block_reg[2][2][9]  ( .D(n2418), .CK(clk), .RN(n3695), .Q(
        \block[2][2][9] ), .QN(n417) );
  DFFRX1 \block_reg[2][2][8]  ( .D(n2419), .CK(clk), .RN(n3695), .Q(
        \block[2][2][8] ), .QN(n416) );
  DFFRX1 \block_reg[2][2][7]  ( .D(n2420), .CK(clk), .RN(n3695), .Q(
        \block[2][2][7] ), .QN(n415) );
  DFFRX1 \block_reg[2][2][6]  ( .D(n2421), .CK(clk), .RN(n3695), .Q(
        \block[2][2][6] ), .QN(n414) );
  DFFRX1 \block_reg[2][2][5]  ( .D(n2422), .CK(clk), .RN(n3695), .Q(
        \block[2][2][5] ), .QN(n413) );
  DFFRX1 \block_reg[2][2][4]  ( .D(n2423), .CK(clk), .RN(n3695), .Q(
        \block[2][2][4] ), .QN(n412) );
  DFFRX1 \block_reg[2][2][3]  ( .D(n2424), .CK(clk), .RN(n3695), .Q(
        \block[2][2][3] ), .QN(n411) );
  DFFRX1 \block_reg[2][2][2]  ( .D(n2425), .CK(clk), .RN(n3695), .Q(
        \block[2][2][2] ), .QN(n410) );
  DFFRX1 \block_reg[2][2][1]  ( .D(n2426), .CK(clk), .RN(n3695), .Q(
        \block[2][2][1] ), .QN(n409) );
  DFFRX1 \block_reg[2][2][0]  ( .D(n2427), .CK(clk), .RN(n3695), .Q(
        \block[2][2][0] ), .QN(n408) );
  DFFRX1 \block_reg[6][1][31]  ( .D(n1916), .CK(clk), .RN(n3687), .Q(
        \block[6][1][31] ), .QN(n919) );
  DFFRX1 \block_reg[6][1][30]  ( .D(n1917), .CK(clk), .RN(n3687), .Q(
        \block[6][1][30] ), .QN(n918) );
  DFFRX1 \block_reg[6][1][29]  ( .D(n1918), .CK(clk), .RN(n3686), .Q(
        \block[6][1][29] ), .QN(n917) );
  DFFRX1 \block_reg[6][1][28]  ( .D(n1919), .CK(clk), .RN(n3686), .Q(
        \block[6][1][28] ), .QN(n916) );
  DFFRX1 \block_reg[6][1][27]  ( .D(n1920), .CK(clk), .RN(n3686), .Q(
        \block[6][1][27] ), .QN(n915) );
  DFFRX1 \block_reg[6][1][26]  ( .D(n1921), .CK(clk), .RN(n3686), .Q(
        \block[6][1][26] ), .QN(n914) );
  DFFRX1 \block_reg[6][1][25]  ( .D(n1922), .CK(clk), .RN(n3686), .Q(
        \block[6][1][25] ), .QN(n913) );
  DFFRX1 \block_reg[6][1][24]  ( .D(n1923), .CK(clk), .RN(n3686), .Q(
        \block[6][1][24] ), .QN(n912) );
  DFFRX1 \block_reg[6][1][23]  ( .D(n1924), .CK(clk), .RN(n3686), .Q(
        \block[6][1][23] ), .QN(n911) );
  DFFRX1 \block_reg[6][1][22]  ( .D(n1925), .CK(clk), .RN(n3686), .Q(
        \block[6][1][22] ), .QN(n910) );
  DFFRX1 \block_reg[6][1][21]  ( .D(n1926), .CK(clk), .RN(n3686), .Q(
        \block[6][1][21] ), .QN(n909) );
  DFFRX1 \block_reg[6][1][20]  ( .D(n1927), .CK(clk), .RN(n3686), .Q(
        \block[6][1][20] ), .QN(n908) );
  DFFRX1 \block_reg[6][1][19]  ( .D(n1928), .CK(clk), .RN(n3686), .Q(
        \block[6][1][19] ), .QN(n907) );
  DFFRX1 \block_reg[6][1][18]  ( .D(n1929), .CK(clk), .RN(n3686), .Q(
        \block[6][1][18] ), .QN(n906) );
  DFFRX1 \block_reg[6][1][17]  ( .D(n1930), .CK(clk), .RN(n3685), .Q(
        \block[6][1][17] ), .QN(n905) );
  DFFRX1 \block_reg[6][1][16]  ( .D(n1931), .CK(clk), .RN(n3685), .Q(
        \block[6][1][16] ), .QN(n904) );
  DFFRX1 \block_reg[6][1][15]  ( .D(n1932), .CK(clk), .RN(n3685), .Q(
        \block[6][1][15] ), .QN(n903) );
  DFFRX1 \block_reg[6][1][14]  ( .D(n1933), .CK(clk), .RN(n3685), .Q(
        \block[6][1][14] ), .QN(n902) );
  DFFRX1 \block_reg[6][1][13]  ( .D(n1934), .CK(clk), .RN(n3685), .Q(
        \block[6][1][13] ), .QN(n901) );
  DFFRX1 \block_reg[6][1][12]  ( .D(n1935), .CK(clk), .RN(n3685), .Q(
        \block[6][1][12] ), .QN(n900) );
  DFFRX1 \block_reg[6][1][11]  ( .D(n1936), .CK(clk), .RN(n3685), .Q(
        \block[6][1][11] ), .QN(n899) );
  DFFRX1 \block_reg[6][1][10]  ( .D(n1937), .CK(clk), .RN(n3685), .Q(
        \block[6][1][10] ), .QN(n898) );
  DFFRX1 \block_reg[6][1][9]  ( .D(n1938), .CK(clk), .RN(n3685), .Q(
        \block[6][1][9] ), .QN(n897) );
  DFFRX1 \block_reg[6][1][8]  ( .D(n1939), .CK(clk), .RN(n3685), .Q(
        \block[6][1][8] ), .QN(n896) );
  DFFRX1 \block_reg[6][1][7]  ( .D(n1940), .CK(clk), .RN(n3685), .Q(
        \block[6][1][7] ), .QN(n895) );
  DFFRX1 \block_reg[6][1][6]  ( .D(n1941), .CK(clk), .RN(n3685), .Q(
        \block[6][1][6] ), .QN(n894) );
  DFFRX1 \block_reg[6][1][5]  ( .D(n1942), .CK(clk), .RN(n3684), .Q(
        \block[6][1][5] ), .QN(n893) );
  DFFRX1 \block_reg[6][1][4]  ( .D(n1943), .CK(clk), .RN(n3684), .Q(
        \block[6][1][4] ), .QN(n892) );
  DFFRX1 \block_reg[6][1][3]  ( .D(n1944), .CK(clk), .RN(n3684), .Q(
        \block[6][1][3] ), .QN(n891) );
  DFFRX1 \block_reg[6][1][2]  ( .D(n1945), .CK(clk), .RN(n3684), .Q(
        \block[6][1][2] ), .QN(n890) );
  DFFRX1 \block_reg[6][1][1]  ( .D(n1946), .CK(clk), .RN(n3684), .Q(
        \block[6][1][1] ), .QN(n889) );
  DFFRX1 \block_reg[6][1][0]  ( .D(n1947), .CK(clk), .RN(n3684), .Q(
        \block[6][1][0] ), .QN(n888) );
  DFFRX1 \block_reg[2][1][24]  ( .D(n2435), .CK(clk), .RN(n3676), .Q(
        \block[2][1][24] ), .QN(n1695) );
  DFFRX1 \block_reg[2][1][23]  ( .D(n2436), .CK(clk), .RN(n3676), .Q(
        \block[2][1][23] ), .QN(n1694) );
  DFFRX1 \block_reg[2][1][22]  ( .D(n2437), .CK(clk), .RN(n3676), .Q(
        \block[2][1][22] ), .QN(n1693) );
  DFFRX1 \block_reg[2][1][21]  ( .D(n2438), .CK(clk), .RN(n3676), .Q(
        \block[2][1][21] ), .QN(n1692) );
  DFFRX1 \block_reg[2][1][20]  ( .D(n2439), .CK(clk), .RN(n3676), .Q(
        \block[2][1][20] ), .QN(n1691) );
  DFFRX1 \block_reg[2][1][19]  ( .D(n2440), .CK(clk), .RN(n3676), .Q(
        \block[2][1][19] ), .QN(n1690) );
  DFFRX1 \block_reg[2][1][18]  ( .D(n2441), .CK(clk), .RN(n3675), .Q(
        \block[2][1][18] ), .QN(n1689) );
  DFFRX1 \block_reg[2][1][17]  ( .D(n2442), .CK(clk), .RN(n3675), .Q(
        \block[2][1][17] ), .QN(n1688) );
  DFFRX1 \block_reg[2][1][16]  ( .D(n2443), .CK(clk), .RN(n3675), .Q(
        \block[2][1][16] ), .QN(n1687) );
  DFFRX1 \block_reg[2][1][15]  ( .D(n2444), .CK(clk), .RN(n3675), .Q(
        \block[2][1][15] ), .QN(n1686) );
  DFFRX1 \block_reg[2][1][14]  ( .D(n2445), .CK(clk), .RN(n3675), .Q(
        \block[2][1][14] ), .QN(n1685) );
  DFFRX1 \block_reg[2][1][13]  ( .D(n2446), .CK(clk), .RN(n3675), .Q(
        \block[2][1][13] ), .QN(n1684) );
  DFFRX1 \block_reg[2][1][12]  ( .D(n2447), .CK(clk), .RN(n3675), .Q(
        \block[2][1][12] ), .QN(n1683) );
  DFFRX1 \block_reg[2][1][11]  ( .D(n2448), .CK(clk), .RN(n3675), .Q(
        \block[2][1][11] ), .QN(n1682) );
  DFFRX1 \block_reg[2][1][10]  ( .D(n2449), .CK(clk), .RN(n3675), .Q(
        \block[2][1][10] ), .QN(n1681) );
  DFFRX1 \block_reg[2][1][9]  ( .D(n2450), .CK(clk), .RN(n3675), .Q(
        \block[2][1][9] ), .QN(n1680) );
  DFFRX1 \block_reg[2][1][8]  ( .D(n2451), .CK(clk), .RN(n3675), .Q(
        \block[2][1][8] ), .QN(n1679) );
  DFFRX1 \block_reg[2][1][7]  ( .D(n2452), .CK(clk), .RN(n3675), .Q(
        \block[2][1][7] ), .QN(n1678) );
  DFFRX1 \block_reg[2][1][6]  ( .D(n2453), .CK(clk), .RN(n3674), .Q(
        \block[2][1][6] ), .QN(n1677) );
  DFFRX1 \block_reg[2][1][5]  ( .D(n2454), .CK(clk), .RN(n3674), .Q(
        \block[2][1][5] ), .QN(n1676) );
  DFFRX1 \block_reg[2][1][4]  ( .D(n2455), .CK(clk), .RN(n3674), .Q(
        \block[2][1][4] ), .QN(n1675) );
  DFFRX1 \block_reg[2][1][3]  ( .D(n2456), .CK(clk), .RN(n3674), .Q(
        \block[2][1][3] ), .QN(n1674) );
  DFFRX1 \block_reg[2][1][2]  ( .D(n2457), .CK(clk), .RN(n3674), .Q(
        \block[2][1][2] ), .QN(n1673) );
  DFFRX1 \block_reg[2][1][1]  ( .D(n2458), .CK(clk), .RN(n3674), .Q(
        \block[2][1][1] ), .QN(n1672) );
  DFFRX1 \block_reg[2][1][0]  ( .D(n2459), .CK(clk), .RN(n3674), .Q(
        \block[2][1][0] ), .QN(n1671) );
  DFFRX1 \block_reg[2][1][31]  ( .D(n2428), .CK(clk), .RN(n3674), .Q(
        \block[2][1][31] ), .QN(n407) );
  DFFRX1 \block_reg[2][1][30]  ( .D(n2429), .CK(clk), .RN(n3674), .Q(
        \block[2][1][30] ), .QN(n406) );
  DFFRX1 \block_reg[2][1][29]  ( .D(n2430), .CK(clk), .RN(n3674), .Q(
        \block[2][1][29] ), .QN(n405) );
  DFFRX1 \block_reg[2][1][28]  ( .D(n2431), .CK(clk), .RN(n3674), .Q(
        \block[2][1][28] ), .QN(n404) );
  DFFRX1 \block_reg[2][1][27]  ( .D(n2432), .CK(clk), .RN(n3674), .Q(
        \block[2][1][27] ), .QN(n403) );
  DFFRX1 \block_reg[2][1][26]  ( .D(n2433), .CK(clk), .RN(n3673), .Q(
        \block[2][1][26] ), .QN(n402) );
  DFFRX1 \block_reg[2][1][25]  ( .D(n2434), .CK(clk), .RN(n3673), .Q(
        \block[2][1][25] ), .QN(n401) );
  DFFRX1 \dirty_reg[7]  ( .D(n1716), .CK(clk), .RN(n3759), .Q(dirty[7]), .QN(
        n1119) );
  DFFRX1 \dirty_reg[3]  ( .D(n1720), .CK(clk), .RN(n3759), .Q(dirty[3]), .QN(
        n1115) );
  DFFRX1 \dirty_reg[5]  ( .D(n1718), .CK(clk), .RN(n3759), .Q(dirty[5]), .QN(
        n1117) );
  DFFRX1 \dirty_reg[1]  ( .D(n1722), .CK(clk), .RN(n3759), .Q(dirty[1]), .QN(
        n1113) );
  DFFRX1 \block_reg[1][0][31]  ( .D(n2588), .CK(clk), .RN(n3756), .Q(
        \block[1][0][31] ), .QN(n1542) );
  DFFRX1 \block_reg[1][0][30]  ( .D(n2589), .CK(clk), .RN(n3756), .Q(
        \block[1][0][30] ), .QN(n1541) );
  DFFRX1 \block_reg[1][0][29]  ( .D(n2590), .CK(clk), .RN(n3756), .Q(
        \block[1][0][29] ), .QN(n1540) );
  DFFRX1 \block_reg[1][0][28]  ( .D(n2591), .CK(clk), .RN(n3756), .Q(
        \block[1][0][28] ), .QN(n1539) );
  DFFRX1 \block_reg[1][0][27]  ( .D(n2592), .CK(clk), .RN(n3756), .Q(
        \block[1][0][27] ), .QN(n1538) );
  DFFRX1 \block_reg[1][0][26]  ( .D(n2593), .CK(clk), .RN(n3756), .Q(
        \block[1][0][26] ), .QN(n1537) );
  DFFRX1 \block_reg[1][0][25]  ( .D(n2594), .CK(clk), .RN(n3755), .Q(
        \block[1][0][25] ), .QN(n1536) );
  DFFRX1 \block_reg[1][0][24]  ( .D(n2595), .CK(clk), .RN(n3755), .Q(
        \block[1][0][24] ), .QN(n1535) );
  DFFRX1 \block_reg[1][0][23]  ( .D(n2596), .CK(clk), .RN(n3755), .Q(
        \block[1][0][23] ), .QN(n1534) );
  DFFRX1 \block_reg[1][0][22]  ( .D(n2597), .CK(clk), .RN(n3755), .Q(
        \block[1][0][22] ), .QN(n1533) );
  DFFRX1 \block_reg[1][0][21]  ( .D(n2598), .CK(clk), .RN(n3755), .Q(
        \block[1][0][21] ), .QN(n1532) );
  DFFRX1 \block_reg[1][0][20]  ( .D(n2599), .CK(clk), .RN(n3755), .Q(
        \block[1][0][20] ), .QN(n1531) );
  DFFRX1 \block_reg[1][0][19]  ( .D(n2600), .CK(clk), .RN(n3755), .Q(
        \block[1][0][19] ), .QN(n1530) );
  DFFRX1 \block_reg[1][0][18]  ( .D(n2601), .CK(clk), .RN(n3755), .Q(
        \block[1][0][18] ), .QN(n1529) );
  DFFRX1 \block_reg[1][0][17]  ( .D(n2602), .CK(clk), .RN(n3755), .Q(
        \block[1][0][17] ), .QN(n1528) );
  DFFRX1 \block_reg[1][0][16]  ( .D(n2603), .CK(clk), .RN(n3755), .Q(
        \block[1][0][16] ), .QN(n1527) );
  DFFRX1 \block_reg[1][0][15]  ( .D(n2604), .CK(clk), .RN(n3755), .Q(
        \block[1][0][15] ), .QN(n1526) );
  DFFRX1 \block_reg[1][0][14]  ( .D(n2605), .CK(clk), .RN(n3755), .Q(
        \block[1][0][14] ), .QN(n1525) );
  DFFRX1 \block_reg[1][0][13]  ( .D(n2606), .CK(clk), .RN(n3754), .Q(
        \block[1][0][13] ), .QN(n1524) );
  DFFRX1 \block_reg[1][0][12]  ( .D(n2607), .CK(clk), .RN(n3754), .Q(
        \block[1][0][12] ), .QN(n1523) );
  DFFRX1 \block_reg[1][0][11]  ( .D(n2608), .CK(clk), .RN(n3754), .Q(
        \block[1][0][11] ), .QN(n1522) );
  DFFRX1 \block_reg[1][0][10]  ( .D(n2609), .CK(clk), .RN(n3754), .Q(
        \block[1][0][10] ), .QN(n1521) );
  DFFRX1 \block_reg[1][0][9]  ( .D(n2610), .CK(clk), .RN(n3754), .Q(
        \block[1][0][9] ), .QN(n1520) );
  DFFRX1 \block_reg[1][0][8]  ( .D(n2611), .CK(clk), .RN(n3754), .Q(
        \block[1][0][8] ), .QN(n1519) );
  DFFRX1 \block_reg[1][0][7]  ( .D(n2612), .CK(clk), .RN(n3754), .Q(
        \block[1][0][7] ), .QN(n1518) );
  DFFRX1 \block_reg[1][0][6]  ( .D(n2613), .CK(clk), .RN(n3754), .Q(
        \block[1][0][6] ), .QN(n1517) );
  DFFRX1 \block_reg[1][0][5]  ( .D(n2614), .CK(clk), .RN(n3754), .Q(
        \block[1][0][5] ), .QN(n1516) );
  DFFRX1 \block_reg[1][0][4]  ( .D(n2615), .CK(clk), .RN(n3754), .Q(
        \block[1][0][4] ), .QN(n1515) );
  DFFRX1 \block_reg[1][0][3]  ( .D(n2616), .CK(clk), .RN(n3754), .Q(
        \block[1][0][3] ), .QN(n1514) );
  DFFRX1 \block_reg[1][0][2]  ( .D(n2617), .CK(clk), .RN(n3754), .Q(
        \block[1][0][2] ), .QN(n1513) );
  DFFRX1 \block_reg[1][0][1]  ( .D(n2618), .CK(clk), .RN(n3753), .Q(
        \block[1][0][1] ), .QN(n1512) );
  DFFRX1 \block_reg[1][0][0]  ( .D(n2619), .CK(clk), .RN(n3753), .Q(
        \block[1][0][0] ), .QN(n1511) );
  DFFRX1 \block_reg[5][0][31]  ( .D(n2076), .CK(clk), .RN(n3745), .Q(
        \block[5][0][31] ), .QN(n759) );
  DFFRX1 \block_reg[5][0][30]  ( .D(n2077), .CK(clk), .RN(n3745), .Q(
        \block[5][0][30] ), .QN(n758) );
  DFFRX1 \block_reg[5][0][29]  ( .D(n2078), .CK(clk), .RN(n3745), .Q(
        \block[5][0][29] ), .QN(n757) );
  DFFRX1 \block_reg[5][0][28]  ( .D(n2079), .CK(clk), .RN(n3745), .Q(
        \block[5][0][28] ), .QN(n756) );
  DFFRX1 \block_reg[5][0][27]  ( .D(n2080), .CK(clk), .RN(n3745), .Q(
        \block[5][0][27] ), .QN(n755) );
  DFFRX1 \block_reg[5][0][26]  ( .D(n2081), .CK(clk), .RN(n3745), .Q(
        \block[5][0][26] ), .QN(n754) );
  DFFRX1 \block_reg[5][0][25]  ( .D(n2082), .CK(clk), .RN(n3745), .Q(
        \block[5][0][25] ), .QN(n753) );
  DFFRX1 \block_reg[5][0][24]  ( .D(n2083), .CK(clk), .RN(n3745), .Q(
        \block[5][0][24] ), .QN(n752) );
  DFFRX1 \block_reg[5][0][23]  ( .D(n2084), .CK(clk), .RN(n3745), .Q(
        \block[5][0][23] ), .QN(n751) );
  DFFRX1 \block_reg[5][0][22]  ( .D(n2085), .CK(clk), .RN(n3745), .Q(
        \block[5][0][22] ), .QN(n750) );
  DFFRX1 \block_reg[5][0][21]  ( .D(n2086), .CK(clk), .RN(n3744), .Q(
        \block[5][0][21] ), .QN(n749) );
  DFFRX1 \block_reg[5][0][20]  ( .D(n2087), .CK(clk), .RN(n3744), .Q(
        \block[5][0][20] ), .QN(n748) );
  DFFRX1 \block_reg[5][0][19]  ( .D(n2088), .CK(clk), .RN(n3744), .Q(
        \block[5][0][19] ), .QN(n747) );
  DFFRX1 \block_reg[5][0][18]  ( .D(n2089), .CK(clk), .RN(n3744), .Q(
        \block[5][0][18] ), .QN(n746) );
  DFFRX1 \block_reg[5][0][17]  ( .D(n2090), .CK(clk), .RN(n3744), .Q(
        \block[5][0][17] ), .QN(n745) );
  DFFRX1 \block_reg[5][0][16]  ( .D(n2091), .CK(clk), .RN(n3744), .Q(
        \block[5][0][16] ), .QN(n744) );
  DFFRX1 \block_reg[5][0][15]  ( .D(n2092), .CK(clk), .RN(n3744), .Q(
        \block[5][0][15] ), .QN(n743) );
  DFFRX1 \block_reg[5][0][14]  ( .D(n2093), .CK(clk), .RN(n3744), .Q(
        \block[5][0][14] ), .QN(n742) );
  DFFRX1 \block_reg[5][0][13]  ( .D(n2094), .CK(clk), .RN(n3744), .Q(
        \block[5][0][13] ), .QN(n741) );
  DFFRX1 \block_reg[5][0][12]  ( .D(n2095), .CK(clk), .RN(n3744), .Q(
        \block[5][0][12] ), .QN(n740) );
  DFFRX1 \block_reg[5][0][11]  ( .D(n2096), .CK(clk), .RN(n3744), .Q(
        \block[5][0][11] ), .QN(n739) );
  DFFRX1 \block_reg[5][0][10]  ( .D(n2097), .CK(clk), .RN(n3744), .Q(
        \block[5][0][10] ), .QN(n738) );
  DFFRX1 \block_reg[5][0][9]  ( .D(n2098), .CK(clk), .RN(n3743), .Q(
        \block[5][0][9] ), .QN(n737) );
  DFFRX1 \block_reg[5][0][8]  ( .D(n2099), .CK(clk), .RN(n3743), .Q(
        \block[5][0][8] ), .QN(n736) );
  DFFRX1 \block_reg[5][0][7]  ( .D(n2100), .CK(clk), .RN(n3743), .Q(
        \block[5][0][7] ), .QN(n735) );
  DFFRX1 \block_reg[5][0][6]  ( .D(n2101), .CK(clk), .RN(n3743), .Q(
        \block[5][0][6] ), .QN(n734) );
  DFFRX1 \block_reg[5][0][5]  ( .D(n2102), .CK(clk), .RN(n3743), .Q(
        \block[5][0][5] ), .QN(n733) );
  DFFRX1 \block_reg[5][0][4]  ( .D(n2103), .CK(clk), .RN(n3743), .Q(
        \block[5][0][4] ), .QN(n732) );
  DFFRX1 \block_reg[5][0][3]  ( .D(n2104), .CK(clk), .RN(n3743), .Q(
        \block[5][0][3] ), .QN(n731) );
  DFFRX1 \block_reg[5][0][2]  ( .D(n2105), .CK(clk), .RN(n3743), .Q(
        \block[5][0][2] ), .QN(n730) );
  DFFRX1 \block_reg[5][0][1]  ( .D(n2106), .CK(clk), .RN(n3743), .Q(
        \block[5][0][1] ), .QN(n729) );
  DFFRX1 \block_reg[5][0][0]  ( .D(n2107), .CK(clk), .RN(n3743), .Q(
        \block[5][0][0] ), .QN(n728) );
  DFFRX1 \block_reg[1][3][31]  ( .D(n2492), .CK(clk), .RN(n3737), .Q(
        \block[1][3][31] ), .QN(n1638) );
  DFFRX1 \block_reg[1][3][30]  ( .D(n2493), .CK(clk), .RN(n3737), .Q(
        \block[1][3][30] ), .QN(n1637) );
  DFFRX1 \block_reg[1][3][29]  ( .D(n2494), .CK(clk), .RN(n3737), .Q(
        \block[1][3][29] ), .QN(n1636) );
  DFFRX1 \block_reg[1][3][28]  ( .D(n2495), .CK(clk), .RN(n3737), .Q(
        \block[1][3][28] ), .QN(n1635) );
  DFFRX1 \block_reg[1][3][27]  ( .D(n2496), .CK(clk), .RN(n3737), .Q(
        \block[1][3][27] ), .QN(n1634) );
  DFFRX1 \block_reg[1][3][26]  ( .D(n2497), .CK(clk), .RN(n3737), .Q(
        \block[1][3][26] ), .QN(n1633) );
  DFFRX1 \block_reg[1][3][25]  ( .D(n2498), .CK(clk), .RN(n3737), .Q(
        \block[1][3][25] ), .QN(n1632) );
  DFFRX1 \block_reg[1][3][24]  ( .D(n2499), .CK(clk), .RN(n3737), .Q(
        \block[1][3][24] ), .QN(n1631) );
  DFFRX1 \block_reg[1][3][23]  ( .D(n2500), .CK(clk), .RN(n3737), .Q(
        \block[1][3][23] ), .QN(n1630) );
  DFFRX1 \block_reg[1][3][22]  ( .D(n2501), .CK(clk), .RN(n3737), .Q(
        \block[1][3][22] ), .QN(n1629) );
  DFFRX1 \block_reg[1][3][21]  ( .D(n2502), .CK(clk), .RN(n3736), .Q(
        \block[1][3][21] ), .QN(n1628) );
  DFFRX1 \block_reg[1][3][20]  ( .D(n2503), .CK(clk), .RN(n3736), .Q(
        \block[1][3][20] ), .QN(n1627) );
  DFFRX1 \block_reg[1][3][19]  ( .D(n2504), .CK(clk), .RN(n3736), .Q(
        \block[1][3][19] ), .QN(n1626) );
  DFFRX1 \block_reg[1][3][18]  ( .D(n2505), .CK(clk), .RN(n3736), .Q(
        \block[1][3][18] ), .QN(n1625) );
  DFFRX1 \block_reg[1][3][17]  ( .D(n2506), .CK(clk), .RN(n3736), .Q(
        \block[1][3][17] ), .QN(n1624) );
  DFFRX1 \block_reg[1][3][16]  ( .D(n2507), .CK(clk), .RN(n3736), .Q(
        \block[1][3][16] ), .QN(n1623) );
  DFFRX1 \block_reg[1][3][15]  ( .D(n2508), .CK(clk), .RN(n3736), .Q(
        \block[1][3][15] ), .QN(n1622) );
  DFFRX1 \block_reg[1][3][14]  ( .D(n2509), .CK(clk), .RN(n3736), .Q(
        \block[1][3][14] ), .QN(n1621) );
  DFFRX1 \block_reg[1][3][13]  ( .D(n2510), .CK(clk), .RN(n3736), .Q(
        \block[1][3][13] ), .QN(n1620) );
  DFFRX1 \block_reg[1][3][12]  ( .D(n2511), .CK(clk), .RN(n3736), .Q(
        \block[1][3][12] ), .QN(n1619) );
  DFFRX1 \block_reg[1][3][11]  ( .D(n2512), .CK(clk), .RN(n3736), .Q(
        \block[1][3][11] ), .QN(n1618) );
  DFFRX1 \block_reg[1][3][10]  ( .D(n2513), .CK(clk), .RN(n3736), .Q(
        \block[1][3][10] ), .QN(n1617) );
  DFFRX1 \block_reg[1][3][9]  ( .D(n2514), .CK(clk), .RN(n3735), .Q(
        \block[1][3][9] ), .QN(n1616) );
  DFFRX1 \block_reg[1][3][8]  ( .D(n2515), .CK(clk), .RN(n3735), .Q(
        \block[1][3][8] ), .QN(n1615) );
  DFFRX1 \block_reg[1][3][7]  ( .D(n2516), .CK(clk), .RN(n3735), .Q(
        \block[1][3][7] ), .QN(n1614) );
  DFFRX1 \block_reg[1][3][6]  ( .D(n2517), .CK(clk), .RN(n3735), .Q(
        \block[1][3][6] ), .QN(n1613) );
  DFFRX1 \block_reg[1][3][5]  ( .D(n2518), .CK(clk), .RN(n3735), .Q(
        \block[1][3][5] ), .QN(n1612) );
  DFFRX1 \block_reg[1][3][4]  ( .D(n2519), .CK(clk), .RN(n3735), .Q(
        \block[1][3][4] ), .QN(n1611) );
  DFFRX1 \block_reg[1][3][3]  ( .D(n2520), .CK(clk), .RN(n3735), .Q(
        \block[1][3][3] ), .QN(n1610) );
  DFFRX1 \block_reg[1][3][2]  ( .D(n2521), .CK(clk), .RN(n3735), .Q(
        \block[1][3][2] ), .QN(n1609) );
  DFFRX1 \block_reg[1][3][1]  ( .D(n2522), .CK(clk), .RN(n3735), .Q(
        \block[1][3][1] ), .QN(n1608) );
  DFFRX1 \block_reg[1][3][0]  ( .D(n2523), .CK(clk), .RN(n3735), .Q(
        \block[1][3][0] ), .QN(n1607) );
  DFFRX1 \block_reg[5][3][31]  ( .D(n1980), .CK(clk), .RN(n3727), .Q(
        \block[5][3][31] ), .QN(n855) );
  DFFRX1 \block_reg[5][3][30]  ( .D(n1981), .CK(clk), .RN(n3727), .Q(
        \block[5][3][30] ), .QN(n854) );
  DFFRX1 \block_reg[5][3][29]  ( .D(n1982), .CK(clk), .RN(n3726), .Q(
        \block[5][3][29] ), .QN(n853) );
  DFFRX1 \block_reg[5][3][28]  ( .D(n1983), .CK(clk), .RN(n3726), .Q(
        \block[5][3][28] ), .QN(n852) );
  DFFRX1 \block_reg[5][3][27]  ( .D(n1984), .CK(clk), .RN(n3726), .Q(
        \block[5][3][27] ), .QN(n851) );
  DFFRX1 \block_reg[5][3][26]  ( .D(n1985), .CK(clk), .RN(n3726), .Q(
        \block[5][3][26] ), .QN(n850) );
  DFFRX1 \block_reg[5][3][25]  ( .D(n1986), .CK(clk), .RN(n3726), .Q(
        \block[5][3][25] ), .QN(n849) );
  DFFRX1 \block_reg[5][3][24]  ( .D(n1987), .CK(clk), .RN(n3726), .Q(
        \block[5][3][24] ), .QN(n848) );
  DFFRX1 \block_reg[5][3][23]  ( .D(n1988), .CK(clk), .RN(n3726), .Q(
        \block[5][3][23] ), .QN(n847) );
  DFFRX1 \block_reg[5][3][22]  ( .D(n1989), .CK(clk), .RN(n3726), .Q(
        \block[5][3][22] ), .QN(n846) );
  DFFRX1 \block_reg[5][3][21]  ( .D(n1990), .CK(clk), .RN(n3726), .Q(
        \block[5][3][21] ), .QN(n845) );
  DFFRX1 \block_reg[5][3][20]  ( .D(n1991), .CK(clk), .RN(n3726), .Q(
        \block[5][3][20] ), .QN(n844) );
  DFFRX1 \block_reg[5][3][19]  ( .D(n1992), .CK(clk), .RN(n3726), .Q(
        \block[5][3][19] ), .QN(n843) );
  DFFRX1 \block_reg[5][3][18]  ( .D(n1993), .CK(clk), .RN(n3726), .Q(
        \block[5][3][18] ), .QN(n842) );
  DFFRX1 \block_reg[5][3][17]  ( .D(n1994), .CK(clk), .RN(n3725), .Q(
        \block[5][3][17] ), .QN(n841) );
  DFFRX1 \block_reg[5][3][16]  ( .D(n1995), .CK(clk), .RN(n3725), .Q(
        \block[5][3][16] ), .QN(n840) );
  DFFRX1 \block_reg[5][3][15]  ( .D(n1996), .CK(clk), .RN(n3725), .Q(
        \block[5][3][15] ), .QN(n839) );
  DFFRX1 \block_reg[5][3][14]  ( .D(n1997), .CK(clk), .RN(n3725), .Q(
        \block[5][3][14] ), .QN(n838) );
  DFFRX1 \block_reg[5][3][13]  ( .D(n1998), .CK(clk), .RN(n3725), .Q(
        \block[5][3][13] ), .QN(n837) );
  DFFRX1 \block_reg[5][3][12]  ( .D(n1999), .CK(clk), .RN(n3725), .Q(
        \block[5][3][12] ), .QN(n836) );
  DFFRX1 \block_reg[5][3][11]  ( .D(n2000), .CK(clk), .RN(n3725), .Q(
        \block[5][3][11] ), .QN(n835) );
  DFFRX1 \block_reg[5][3][10]  ( .D(n2001), .CK(clk), .RN(n3725), .Q(
        \block[5][3][10] ), .QN(n834) );
  DFFRX1 \block_reg[5][3][9]  ( .D(n2002), .CK(clk), .RN(n3725), .Q(
        \block[5][3][9] ), .QN(n833) );
  DFFRX1 \block_reg[5][3][8]  ( .D(n2003), .CK(clk), .RN(n3725), .Q(
        \block[5][3][8] ), .QN(n832) );
  DFFRX1 \block_reg[5][3][7]  ( .D(n2004), .CK(clk), .RN(n3725), .Q(
        \block[5][3][7] ), .QN(n831) );
  DFFRX1 \block_reg[5][3][6]  ( .D(n2005), .CK(clk), .RN(n3725), .Q(
        \block[5][3][6] ), .QN(n830) );
  DFFRX1 \block_reg[5][3][5]  ( .D(n2006), .CK(clk), .RN(n3724), .Q(
        \block[5][3][5] ), .QN(n829) );
  DFFRX1 \block_reg[5][3][4]  ( .D(n2007), .CK(clk), .RN(n3724), .Q(
        \block[5][3][4] ), .QN(n828) );
  DFFRX1 \block_reg[5][3][3]  ( .D(n2008), .CK(clk), .RN(n3724), .Q(
        \block[5][3][3] ), .QN(n827) );
  DFFRX1 \block_reg[5][3][2]  ( .D(n2009), .CK(clk), .RN(n3724), .Q(
        \block[5][3][2] ), .QN(n826) );
  DFFRX1 \block_reg[5][3][1]  ( .D(n2010), .CK(clk), .RN(n3724), .Q(
        \block[5][3][1] ), .QN(n825) );
  DFFRX1 \block_reg[5][3][0]  ( .D(n2011), .CK(clk), .RN(n3724), .Q(
        \block[5][3][0] ), .QN(n824) );
  DFFRX1 \block_reg[1][2][31]  ( .D(n2524), .CK(clk), .RN(n3716), .Q(
        \block[1][2][31] ), .QN(n1606) );
  DFFRX1 \block_reg[1][2][30]  ( .D(n2525), .CK(clk), .RN(n3716), .Q(
        \block[1][2][30] ), .QN(n1605) );
  DFFRX1 \block_reg[1][2][29]  ( .D(n2526), .CK(clk), .RN(n3716), .Q(
        \block[1][2][29] ), .QN(n1604) );
  DFFRX1 \block_reg[1][2][28]  ( .D(n2527), .CK(clk), .RN(n3716), .Q(
        \block[1][2][28] ), .QN(n1603) );
  DFFRX1 \block_reg[1][2][27]  ( .D(n2528), .CK(clk), .RN(n3716), .Q(
        \block[1][2][27] ), .QN(n1602) );
  DFFRX1 \block_reg[1][2][26]  ( .D(n2529), .CK(clk), .RN(n3716), .Q(
        \block[1][2][26] ), .QN(n1601) );
  DFFRX1 \block_reg[1][2][25]  ( .D(n2530), .CK(clk), .RN(n3715), .Q(
        \block[1][2][25] ), .QN(n1600) );
  DFFRX1 \block_reg[1][2][24]  ( .D(n2531), .CK(clk), .RN(n3715), .Q(
        \block[1][2][24] ), .QN(n1599) );
  DFFRX1 \block_reg[1][2][23]  ( .D(n2532), .CK(clk), .RN(n3715), .Q(
        \block[1][2][23] ), .QN(n1598) );
  DFFRX1 \block_reg[1][2][22]  ( .D(n2533), .CK(clk), .RN(n3715), .Q(
        \block[1][2][22] ), .QN(n1597) );
  DFFRX1 \block_reg[1][2][21]  ( .D(n2534), .CK(clk), .RN(n3715), .Q(
        \block[1][2][21] ), .QN(n1596) );
  DFFRX1 \block_reg[1][2][20]  ( .D(n2535), .CK(clk), .RN(n3715), .Q(
        \block[1][2][20] ), .QN(n1595) );
  DFFRX1 \block_reg[1][2][19]  ( .D(n2536), .CK(clk), .RN(n3715), .Q(
        \block[1][2][19] ), .QN(n1594) );
  DFFRX1 \block_reg[1][2][18]  ( .D(n2537), .CK(clk), .RN(n3715), .Q(
        \block[1][2][18] ), .QN(n1593) );
  DFFRX1 \block_reg[1][2][17]  ( .D(n2538), .CK(clk), .RN(n3715), .Q(
        \block[1][2][17] ), .QN(n1592) );
  DFFRX1 \block_reg[1][2][16]  ( .D(n2539), .CK(clk), .RN(n3715), .Q(
        \block[1][2][16] ), .QN(n1591) );
  DFFRX1 \block_reg[1][2][15]  ( .D(n2540), .CK(clk), .RN(n3715), .Q(
        \block[1][2][15] ), .QN(n1590) );
  DFFRX1 \block_reg[1][2][14]  ( .D(n2541), .CK(clk), .RN(n3715), .Q(
        \block[1][2][14] ), .QN(n1589) );
  DFFRX1 \block_reg[1][2][13]  ( .D(n2542), .CK(clk), .RN(n3714), .Q(
        \block[1][2][13] ), .QN(n1588) );
  DFFRX1 \block_reg[1][2][12]  ( .D(n2543), .CK(clk), .RN(n3714), .Q(
        \block[1][2][12] ), .QN(n1587) );
  DFFRX1 \block_reg[1][2][11]  ( .D(n2544), .CK(clk), .RN(n3714), .Q(
        \block[1][2][11] ), .QN(n1586) );
  DFFRX1 \block_reg[1][2][10]  ( .D(n2545), .CK(clk), .RN(n3714), .Q(
        \block[1][2][10] ), .QN(n1585) );
  DFFRX1 \block_reg[1][2][9]  ( .D(n2546), .CK(clk), .RN(n3714), .Q(
        \block[1][2][9] ), .QN(n1584) );
  DFFRX1 \block_reg[1][2][8]  ( .D(n2547), .CK(clk), .RN(n3714), .Q(
        \block[1][2][8] ), .QN(n1583) );
  DFFRX1 \block_reg[1][2][7]  ( .D(n2548), .CK(clk), .RN(n3714), .Q(
        \block[1][2][7] ), .QN(n1582) );
  DFFRX1 \block_reg[1][2][6]  ( .D(n2549), .CK(clk), .RN(n3714), .Q(
        \block[1][2][6] ), .QN(n1581) );
  DFFRX1 \block_reg[1][2][5]  ( .D(n2550), .CK(clk), .RN(n3714), .Q(
        \block[1][2][5] ), .QN(n1580) );
  DFFRX1 \block_reg[1][2][4]  ( .D(n2551), .CK(clk), .RN(n3714), .Q(
        \block[1][2][4] ), .QN(n1579) );
  DFFRX1 \block_reg[1][2][3]  ( .D(n2552), .CK(clk), .RN(n3714), .Q(
        \block[1][2][3] ), .QN(n1578) );
  DFFRX1 \block_reg[1][2][2]  ( .D(n2553), .CK(clk), .RN(n3714), .Q(
        \block[1][2][2] ), .QN(n1577) );
  DFFRX1 \block_reg[1][2][1]  ( .D(n2554), .CK(clk), .RN(n3713), .Q(
        \block[1][2][1] ), .QN(n1576) );
  DFFRX1 \block_reg[1][2][0]  ( .D(n2555), .CK(clk), .RN(n3713), .Q(
        \block[1][2][0] ), .QN(n1575) );
  DFFRX1 \block_reg[5][2][31]  ( .D(n2012), .CK(clk), .RN(n3705), .Q(
        \block[5][2][31] ), .QN(n823) );
  DFFRX1 \block_reg[5][2][30]  ( .D(n2013), .CK(clk), .RN(n3705), .Q(
        \block[5][2][30] ), .QN(n822) );
  DFFRX1 \block_reg[5][2][29]  ( .D(n2014), .CK(clk), .RN(n3705), .Q(
        \block[5][2][29] ), .QN(n821) );
  DFFRX1 \block_reg[5][2][28]  ( .D(n2015), .CK(clk), .RN(n3705), .Q(
        \block[5][2][28] ), .QN(n820) );
  DFFRX1 \block_reg[5][2][27]  ( .D(n2016), .CK(clk), .RN(n3705), .Q(
        \block[5][2][27] ), .QN(n819) );
  DFFRX1 \block_reg[5][2][26]  ( .D(n2017), .CK(clk), .RN(n3705), .Q(
        \block[5][2][26] ), .QN(n818) );
  DFFRX1 \block_reg[5][2][25]  ( .D(n2018), .CK(clk), .RN(n3705), .Q(
        \block[5][2][25] ), .QN(n817) );
  DFFRX1 \block_reg[5][2][24]  ( .D(n2019), .CK(clk), .RN(n3705), .Q(
        \block[5][2][24] ), .QN(n816) );
  DFFRX1 \block_reg[5][2][23]  ( .D(n2020), .CK(clk), .RN(n3705), .Q(
        \block[5][2][23] ), .QN(n815) );
  DFFRX1 \block_reg[5][2][22]  ( .D(n2021), .CK(clk), .RN(n3705), .Q(
        \block[5][2][22] ), .QN(n814) );
  DFFRX1 \block_reg[5][2][21]  ( .D(n2022), .CK(clk), .RN(n3704), .Q(
        \block[5][2][21] ), .QN(n813) );
  DFFRX1 \block_reg[5][2][20]  ( .D(n2023), .CK(clk), .RN(n3704), .Q(
        \block[5][2][20] ), .QN(n812) );
  DFFRX1 \block_reg[5][2][19]  ( .D(n2024), .CK(clk), .RN(n3704), .Q(
        \block[5][2][19] ), .QN(n811) );
  DFFRX1 \block_reg[5][2][18]  ( .D(n2025), .CK(clk), .RN(n3704), .Q(
        \block[5][2][18] ), .QN(n810) );
  DFFRX1 \block_reg[5][2][17]  ( .D(n2026), .CK(clk), .RN(n3704), .Q(
        \block[5][2][17] ), .QN(n809) );
  DFFRX1 \block_reg[5][2][16]  ( .D(n2027), .CK(clk), .RN(n3704), .Q(
        \block[5][2][16] ), .QN(n808) );
  DFFRX1 \block_reg[5][2][15]  ( .D(n2028), .CK(clk), .RN(n3704), .Q(
        \block[5][2][15] ), .QN(n807) );
  DFFRX1 \block_reg[5][2][14]  ( .D(n2029), .CK(clk), .RN(n3704), .Q(
        \block[5][2][14] ), .QN(n806) );
  DFFRX1 \block_reg[5][2][13]  ( .D(n2030), .CK(clk), .RN(n3704), .Q(
        \block[5][2][13] ), .QN(n805) );
  DFFRX1 \block_reg[5][2][12]  ( .D(n2031), .CK(clk), .RN(n3704), .Q(
        \block[5][2][12] ), .QN(n804) );
  DFFRX1 \block_reg[5][2][11]  ( .D(n2032), .CK(clk), .RN(n3704), .Q(
        \block[5][2][11] ), .QN(n803) );
  DFFRX1 \block_reg[5][2][10]  ( .D(n2033), .CK(clk), .RN(n3704), .Q(
        \block[5][2][10] ), .QN(n802) );
  DFFRX1 \block_reg[5][2][9]  ( .D(n2034), .CK(clk), .RN(n3703), .Q(
        \block[5][2][9] ), .QN(n801) );
  DFFRX1 \block_reg[5][2][8]  ( .D(n2035), .CK(clk), .RN(n3703), .Q(
        \block[5][2][8] ), .QN(n800) );
  DFFRX1 \block_reg[5][2][7]  ( .D(n2036), .CK(clk), .RN(n3703), .Q(
        \block[5][2][7] ), .QN(n799) );
  DFFRX1 \block_reg[5][2][6]  ( .D(n2037), .CK(clk), .RN(n3703), .Q(
        \block[5][2][6] ), .QN(n798) );
  DFFRX1 \block_reg[5][2][5]  ( .D(n2038), .CK(clk), .RN(n3703), .Q(
        \block[5][2][5] ), .QN(n797) );
  DFFRX1 \block_reg[5][2][4]  ( .D(n2039), .CK(clk), .RN(n3703), .Q(
        \block[5][2][4] ), .QN(n796) );
  DFFRX1 \block_reg[5][2][3]  ( .D(n2040), .CK(clk), .RN(n3703), .Q(
        \block[5][2][3] ), .QN(n795) );
  DFFRX1 \block_reg[5][2][2]  ( .D(n2041), .CK(clk), .RN(n3703), .Q(
        \block[5][2][2] ), .QN(n794) );
  DFFRX1 \block_reg[5][2][1]  ( .D(n2042), .CK(clk), .RN(n3703), .Q(
        \block[5][2][1] ), .QN(n793) );
  DFFRX1 \block_reg[5][2][0]  ( .D(n2043), .CK(clk), .RN(n3703), .Q(
        \block[5][2][0] ), .QN(n792) );
  DFFRX1 \block_reg[1][1][31]  ( .D(n2556), .CK(clk), .RN(n3695), .Q(
        \block[1][1][31] ), .QN(n1574) );
  DFFRX1 \block_reg[1][1][30]  ( .D(n2557), .CK(clk), .RN(n3695), .Q(
        \block[1][1][30] ), .QN(n1573) );
  DFFRX1 \block_reg[1][1][29]  ( .D(n2558), .CK(clk), .RN(n3694), .Q(
        \block[1][1][29] ), .QN(n1572) );
  DFFRX1 \block_reg[1][1][28]  ( .D(n2559), .CK(clk), .RN(n3694), .Q(
        \block[1][1][28] ), .QN(n1571) );
  DFFRX1 \block_reg[1][1][27]  ( .D(n2560), .CK(clk), .RN(n3694), .Q(
        \block[1][1][27] ), .QN(n1570) );
  DFFRX1 \block_reg[1][1][26]  ( .D(n2561), .CK(clk), .RN(n3694), .Q(
        \block[1][1][26] ), .QN(n1569) );
  DFFRX1 \block_reg[1][1][25]  ( .D(n2562), .CK(clk), .RN(n3694), .Q(
        \block[1][1][25] ), .QN(n1568) );
  DFFRX1 \block_reg[1][1][24]  ( .D(n2563), .CK(clk), .RN(n3694), .Q(
        \block[1][1][24] ), .QN(n1567) );
  DFFRX1 \block_reg[1][1][23]  ( .D(n2564), .CK(clk), .RN(n3694), .Q(
        \block[1][1][23] ), .QN(n1566) );
  DFFRX1 \block_reg[1][1][22]  ( .D(n2565), .CK(clk), .RN(n3694), .Q(
        \block[1][1][22] ), .QN(n1565) );
  DFFRX1 \block_reg[1][1][21]  ( .D(n2566), .CK(clk), .RN(n3694), .Q(
        \block[1][1][21] ), .QN(n1564) );
  DFFRX1 \block_reg[1][1][20]  ( .D(n2567), .CK(clk), .RN(n3694), .Q(
        \block[1][1][20] ), .QN(n1563) );
  DFFRX1 \block_reg[1][1][19]  ( .D(n2568), .CK(clk), .RN(n3694), .Q(
        \block[1][1][19] ), .QN(n1562) );
  DFFRX1 \block_reg[1][1][18]  ( .D(n2569), .CK(clk), .RN(n3694), .Q(
        \block[1][1][18] ), .QN(n1561) );
  DFFRX1 \block_reg[1][1][17]  ( .D(n2570), .CK(clk), .RN(n3693), .Q(
        \block[1][1][17] ), .QN(n1560) );
  DFFRX1 \block_reg[1][1][16]  ( .D(n2571), .CK(clk), .RN(n3693), .Q(
        \block[1][1][16] ), .QN(n1559) );
  DFFRX1 \block_reg[1][1][15]  ( .D(n2572), .CK(clk), .RN(n3693), .Q(
        \block[1][1][15] ), .QN(n1558) );
  DFFRX1 \block_reg[1][1][14]  ( .D(n2573), .CK(clk), .RN(n3693), .Q(
        \block[1][1][14] ), .QN(n1557) );
  DFFRX1 \block_reg[1][1][13]  ( .D(n2574), .CK(clk), .RN(n3693), .Q(
        \block[1][1][13] ), .QN(n1556) );
  DFFRX1 \block_reg[1][1][12]  ( .D(n2575), .CK(clk), .RN(n3693), .Q(
        \block[1][1][12] ), .QN(n1555) );
  DFFRX1 \block_reg[1][1][11]  ( .D(n2576), .CK(clk), .RN(n3693), .Q(
        \block[1][1][11] ), .QN(n1554) );
  DFFRX1 \block_reg[1][1][10]  ( .D(n2577), .CK(clk), .RN(n3693), .Q(
        \block[1][1][10] ), .QN(n1553) );
  DFFRX1 \block_reg[1][1][9]  ( .D(n2578), .CK(clk), .RN(n3693), .Q(
        \block[1][1][9] ), .QN(n1552) );
  DFFRX1 \block_reg[1][1][8]  ( .D(n2579), .CK(clk), .RN(n3693), .Q(
        \block[1][1][8] ), .QN(n1551) );
  DFFRX1 \block_reg[1][1][7]  ( .D(n2580), .CK(clk), .RN(n3693), .Q(
        \block[1][1][7] ), .QN(n1550) );
  DFFRX1 \block_reg[1][1][6]  ( .D(n2581), .CK(clk), .RN(n3693), .Q(
        \block[1][1][6] ), .QN(n1549) );
  DFFRX1 \block_reg[1][1][5]  ( .D(n2582), .CK(clk), .RN(n3692), .Q(
        \block[1][1][5] ), .QN(n1548) );
  DFFRX1 \block_reg[1][1][4]  ( .D(n2583), .CK(clk), .RN(n3692), .Q(
        \block[1][1][4] ), .QN(n1547) );
  DFFRX1 \block_reg[1][1][3]  ( .D(n2584), .CK(clk), .RN(n3692), .Q(
        \block[1][1][3] ), .QN(n1546) );
  DFFRX1 \block_reg[1][1][2]  ( .D(n2585), .CK(clk), .RN(n3692), .Q(
        \block[1][1][2] ), .QN(n1545) );
  DFFRX1 \block_reg[1][1][1]  ( .D(n2586), .CK(clk), .RN(n3692), .Q(
        \block[1][1][1] ), .QN(n1544) );
  DFFRX1 \block_reg[1][1][0]  ( .D(n2587), .CK(clk), .RN(n3692), .Q(
        \block[1][1][0] ), .QN(n1543) );
  DFFRX1 \block_reg[5][1][31]  ( .D(n2044), .CK(clk), .RN(n3684), .Q(
        \block[5][1][31] ), .QN(n791) );
  DFFRX1 \block_reg[5][1][30]  ( .D(n2045), .CK(clk), .RN(n3684), .Q(
        \block[5][1][30] ), .QN(n790) );
  DFFRX1 \block_reg[5][1][29]  ( .D(n2046), .CK(clk), .RN(n3684), .Q(
        \block[5][1][29] ), .QN(n789) );
  DFFRX1 \block_reg[5][1][28]  ( .D(n2047), .CK(clk), .RN(n3684), .Q(
        \block[5][1][28] ), .QN(n788) );
  DFFRX1 \block_reg[5][1][27]  ( .D(n2048), .CK(clk), .RN(n3684), .Q(
        \block[5][1][27] ), .QN(n787) );
  DFFRX1 \block_reg[5][1][26]  ( .D(n2049), .CK(clk), .RN(n3684), .Q(
        \block[5][1][26] ), .QN(n786) );
  DFFRX1 \block_reg[5][1][25]  ( .D(n2050), .CK(clk), .RN(n3683), .Q(
        \block[5][1][25] ), .QN(n785) );
  DFFRX1 \block_reg[5][1][24]  ( .D(n2051), .CK(clk), .RN(n3683), .Q(
        \block[5][1][24] ), .QN(n784) );
  DFFRX1 \block_reg[5][1][23]  ( .D(n2052), .CK(clk), .RN(n3683), .Q(
        \block[5][1][23] ), .QN(n783) );
  DFFRX1 \block_reg[5][1][22]  ( .D(n2053), .CK(clk), .RN(n3683), .Q(
        \block[5][1][22] ), .QN(n782) );
  DFFRX1 \block_reg[5][1][21]  ( .D(n2054), .CK(clk), .RN(n3683), .Q(
        \block[5][1][21] ), .QN(n781) );
  DFFRX1 \block_reg[5][1][20]  ( .D(n2055), .CK(clk), .RN(n3683), .Q(
        \block[5][1][20] ), .QN(n780) );
  DFFRX1 \block_reg[5][1][19]  ( .D(n2056), .CK(clk), .RN(n3683), .Q(
        \block[5][1][19] ), .QN(n779) );
  DFFRX1 \block_reg[5][1][18]  ( .D(n2057), .CK(clk), .RN(n3683), .Q(
        \block[5][1][18] ), .QN(n778) );
  DFFRX1 \block_reg[5][1][17]  ( .D(n2058), .CK(clk), .RN(n3683), .Q(
        \block[5][1][17] ), .QN(n777) );
  DFFRX1 \block_reg[5][1][16]  ( .D(n2059), .CK(clk), .RN(n3683), .Q(
        \block[5][1][16] ), .QN(n776) );
  DFFRX1 \block_reg[5][1][15]  ( .D(n2060), .CK(clk), .RN(n3683), .Q(
        \block[5][1][15] ), .QN(n775) );
  DFFRX1 \block_reg[5][1][14]  ( .D(n2061), .CK(clk), .RN(n3683), .Q(
        \block[5][1][14] ), .QN(n774) );
  DFFRX1 \block_reg[5][1][13]  ( .D(n2062), .CK(clk), .RN(n3682), .Q(
        \block[5][1][13] ), .QN(n773) );
  DFFRX1 \block_reg[5][1][12]  ( .D(n2063), .CK(clk), .RN(n3682), .Q(
        \block[5][1][12] ), .QN(n772) );
  DFFRX1 \block_reg[5][1][11]  ( .D(n2064), .CK(clk), .RN(n3682), .Q(
        \block[5][1][11] ), .QN(n771) );
  DFFRX1 \block_reg[5][1][10]  ( .D(n2065), .CK(clk), .RN(n3682), .Q(
        \block[5][1][10] ), .QN(n770) );
  DFFRX1 \block_reg[5][1][9]  ( .D(n2066), .CK(clk), .RN(n3682), .Q(
        \block[5][1][9] ), .QN(n769) );
  DFFRX1 \block_reg[5][1][8]  ( .D(n2067), .CK(clk), .RN(n3682), .Q(
        \block[5][1][8] ), .QN(n768) );
  DFFRX1 \block_reg[5][1][7]  ( .D(n2068), .CK(clk), .RN(n3682), .Q(
        \block[5][1][7] ), .QN(n767) );
  DFFRX1 \block_reg[5][1][6]  ( .D(n2069), .CK(clk), .RN(n3682), .Q(
        \block[5][1][6] ), .QN(n766) );
  DFFRX1 \block_reg[5][1][5]  ( .D(n2070), .CK(clk), .RN(n3682), .Q(
        \block[5][1][5] ), .QN(n765) );
  DFFRX1 \block_reg[5][1][4]  ( .D(n2071), .CK(clk), .RN(n3682), .Q(
        \block[5][1][4] ), .QN(n764) );
  DFFRX1 \block_reg[5][1][3]  ( .D(n2072), .CK(clk), .RN(n3682), .Q(
        \block[5][1][3] ), .QN(n763) );
  DFFRX1 \block_reg[5][1][2]  ( .D(n2073), .CK(clk), .RN(n3682), .Q(
        \block[5][1][2] ), .QN(n762) );
  DFFRX1 \block_reg[5][1][1]  ( .D(n2074), .CK(clk), .RN(n3681), .Q(
        \block[5][1][1] ), .QN(n761) );
  DFFRX1 \block_reg[5][1][0]  ( .D(n2075), .CK(clk), .RN(n3681), .Q(
        \block[5][1][0] ), .QN(n760) );
  DFFRX1 \dirty_reg[4]  ( .D(n1719), .CK(clk), .RN(n3759), .Q(dirty[4]), .QN(
        n1116) );
  DFFRX1 \dirty_reg[0]  ( .D(n1723), .CK(clk), .RN(n3759), .Q(dirty[0]), .QN(
        n1112) );
  DFFRX1 \block_reg[0][0][31]  ( .D(n2716), .CK(clk), .RN(n3753), .Q(
        \block[0][0][31] ), .QN(n1414) );
  DFFRX1 \block_reg[0][0][30]  ( .D(n2717), .CK(clk), .RN(n3753), .Q(
        \block[0][0][30] ), .QN(n1413) );
  DFFRX1 \block_reg[0][0][29]  ( .D(n2718), .CK(clk), .RN(n3753), .Q(
        \block[0][0][29] ), .QN(n1412) );
  DFFRX1 \block_reg[0][0][28]  ( .D(n2719), .CK(clk), .RN(n3753), .Q(
        \block[0][0][28] ), .QN(n1411) );
  DFFRX1 \block_reg[0][0][27]  ( .D(n2720), .CK(clk), .RN(n3753), .Q(
        \block[0][0][27] ), .QN(n1410) );
  DFFRX1 \block_reg[0][0][26]  ( .D(n2721), .CK(clk), .RN(n3753), .Q(
        \block[0][0][26] ), .QN(n1409) );
  DFFRX1 \block_reg[0][0][25]  ( .D(n2722), .CK(clk), .RN(n3753), .Q(
        \block[0][0][25] ), .QN(n1408) );
  DFFRX1 \block_reg[0][0][24]  ( .D(n2723), .CK(clk), .RN(n3753), .Q(
        \block[0][0][24] ), .QN(n1407) );
  DFFRX1 \block_reg[0][0][23]  ( .D(n2724), .CK(clk), .RN(n3753), .Q(
        \block[0][0][23] ), .QN(n1406) );
  DFFRX1 \block_reg[0][0][22]  ( .D(n2725), .CK(clk), .RN(n3753), .Q(
        \block[0][0][22] ), .QN(n1405) );
  DFFRX1 \block_reg[0][0][21]  ( .D(n2726), .CK(clk), .RN(n3752), .Q(
        \block[0][0][21] ), .QN(n1404) );
  DFFRX1 \block_reg[0][0][20]  ( .D(n2727), .CK(clk), .RN(n3752), .Q(
        \block[0][0][20] ), .QN(n1403) );
  DFFRX1 \block_reg[0][0][19]  ( .D(n2728), .CK(clk), .RN(n3752), .Q(
        \block[0][0][19] ), .QN(n1402) );
  DFFRX1 \block_reg[0][0][18]  ( .D(n2729), .CK(clk), .RN(n3752), .Q(
        \block[0][0][18] ), .QN(n1401) );
  DFFRX1 \block_reg[0][0][17]  ( .D(n2730), .CK(clk), .RN(n3752), .Q(
        \block[0][0][17] ), .QN(n1400) );
  DFFRX1 \block_reg[0][0][16]  ( .D(n2731), .CK(clk), .RN(n3752), .Q(
        \block[0][0][16] ), .QN(n1399) );
  DFFRX1 \block_reg[0][0][15]  ( .D(n2732), .CK(clk), .RN(n3752), .Q(
        \block[0][0][15] ), .QN(n1398) );
  DFFRX1 \block_reg[0][0][14]  ( .D(n2733), .CK(clk), .RN(n3752), .Q(
        \block[0][0][14] ), .QN(n1397) );
  DFFRX1 \block_reg[0][0][13]  ( .D(n2734), .CK(clk), .RN(n3752), .Q(
        \block[0][0][13] ), .QN(n1396) );
  DFFRX1 \block_reg[0][0][12]  ( .D(n2735), .CK(clk), .RN(n3752), .Q(
        \block[0][0][12] ), .QN(n1395) );
  DFFRX1 \block_reg[0][0][11]  ( .D(n2736), .CK(clk), .RN(n3752), .Q(
        \block[0][0][11] ), .QN(n1394) );
  DFFRX1 \block_reg[0][0][10]  ( .D(n2737), .CK(clk), .RN(n3752), .Q(
        \block[0][0][10] ), .QN(n1393) );
  DFFRX1 \block_reg[0][0][9]  ( .D(n2738), .CK(clk), .RN(n3751), .Q(
        \block[0][0][9] ), .QN(n1392) );
  DFFRX1 \block_reg[0][0][8]  ( .D(n2739), .CK(clk), .RN(n3751), .Q(
        \block[0][0][8] ), .QN(n1391) );
  DFFRX1 \block_reg[0][0][7]  ( .D(n2740), .CK(clk), .RN(n3751), .Q(
        \block[0][0][7] ), .QN(n1390) );
  DFFRX1 \block_reg[0][0][6]  ( .D(n2741), .CK(clk), .RN(n3751), .Q(
        \block[0][0][6] ), .QN(n1389) );
  DFFRX1 \block_reg[0][0][5]  ( .D(n2742), .CK(clk), .RN(n3751), .Q(
        \block[0][0][5] ), .QN(n1388) );
  DFFRX1 \block_reg[0][0][4]  ( .D(n2743), .CK(clk), .RN(n3751), .Q(
        \block[0][0][4] ), .QN(n1387) );
  DFFRX1 \block_reg[0][0][3]  ( .D(n2744), .CK(clk), .RN(n3751), .Q(
        \block[0][0][3] ), .QN(n1386) );
  DFFRX1 \block_reg[0][0][2]  ( .D(n2745), .CK(clk), .RN(n3751), .Q(
        \block[0][0][2] ), .QN(n1385) );
  DFFRX1 \block_reg[0][0][1]  ( .D(n2746), .CK(clk), .RN(n3751), .Q(
        \block[0][0][1] ), .QN(n1384) );
  DFFRX1 \block_reg[0][0][0]  ( .D(n2747), .CK(clk), .RN(n3751), .Q(
        \block[0][0][0] ), .QN(n1383) );
  DFFRX1 \block_reg[4][0][31]  ( .D(n2204), .CK(clk), .RN(n3743), .Q(
        \block[4][0][31] ), .QN(n631) );
  DFFRX1 \block_reg[4][0][30]  ( .D(n2205), .CK(clk), .RN(n3743), .Q(
        \block[4][0][30] ), .QN(n630) );
  DFFRX1 \block_reg[4][0][29]  ( .D(n2206), .CK(clk), .RN(n3742), .Q(
        \block[4][0][29] ), .QN(n629) );
  DFFRX1 \block_reg[4][0][28]  ( .D(n2207), .CK(clk), .RN(n3742), .Q(
        \block[4][0][28] ), .QN(n628) );
  DFFRX1 \block_reg[4][0][27]  ( .D(n2208), .CK(clk), .RN(n3742), .Q(
        \block[4][0][27] ), .QN(n627) );
  DFFRX1 \block_reg[4][0][26]  ( .D(n2209), .CK(clk), .RN(n3742), .Q(
        \block[4][0][26] ), .QN(n626) );
  DFFRX1 \block_reg[4][0][25]  ( .D(n2210), .CK(clk), .RN(n3742), .Q(
        \block[4][0][25] ), .QN(n625) );
  DFFRX1 \block_reg[4][0][24]  ( .D(n2211), .CK(clk), .RN(n3742), .Q(
        \block[4][0][24] ), .QN(n624) );
  DFFRX1 \block_reg[4][0][23]  ( .D(n2212), .CK(clk), .RN(n3742), .Q(
        \block[4][0][23] ), .QN(n623) );
  DFFRX1 \block_reg[4][0][22]  ( .D(n2213), .CK(clk), .RN(n3742), .Q(
        \block[4][0][22] ), .QN(n622) );
  DFFRX1 \block_reg[4][0][21]  ( .D(n2214), .CK(clk), .RN(n3742), .Q(
        \block[4][0][21] ), .QN(n621) );
  DFFRX1 \block_reg[4][0][20]  ( .D(n2215), .CK(clk), .RN(n3742), .Q(
        \block[4][0][20] ), .QN(n620) );
  DFFRX1 \block_reg[4][0][19]  ( .D(n2216), .CK(clk), .RN(n3742), .Q(
        \block[4][0][19] ), .QN(n619) );
  DFFRX1 \block_reg[4][0][18]  ( .D(n2217), .CK(clk), .RN(n3742), .Q(
        \block[4][0][18] ), .QN(n618) );
  DFFRX1 \block_reg[4][0][17]  ( .D(n2218), .CK(clk), .RN(n3741), .Q(
        \block[4][0][17] ), .QN(n617) );
  DFFRX1 \block_reg[4][0][16]  ( .D(n2219), .CK(clk), .RN(n3741), .Q(
        \block[4][0][16] ), .QN(n616) );
  DFFRX1 \block_reg[4][0][15]  ( .D(n2220), .CK(clk), .RN(n3741), .Q(
        \block[4][0][15] ), .QN(n615) );
  DFFRX1 \block_reg[4][0][14]  ( .D(n2221), .CK(clk), .RN(n3741), .Q(
        \block[4][0][14] ), .QN(n614) );
  DFFRX1 \block_reg[4][0][13]  ( .D(n2222), .CK(clk), .RN(n3741), .Q(
        \block[4][0][13] ), .QN(n613) );
  DFFRX1 \block_reg[4][0][12]  ( .D(n2223), .CK(clk), .RN(n3741), .Q(
        \block[4][0][12] ), .QN(n612) );
  DFFRX1 \block_reg[4][0][11]  ( .D(n2224), .CK(clk), .RN(n3741), .Q(
        \block[4][0][11] ), .QN(n611) );
  DFFRX1 \block_reg[4][0][10]  ( .D(n2225), .CK(clk), .RN(n3741), .Q(
        \block[4][0][10] ), .QN(n610) );
  DFFRX1 \block_reg[4][0][9]  ( .D(n2226), .CK(clk), .RN(n3741), .Q(
        \block[4][0][9] ), .QN(n609) );
  DFFRX1 \block_reg[4][0][8]  ( .D(n2227), .CK(clk), .RN(n3741), .Q(
        \block[4][0][8] ), .QN(n608) );
  DFFRX1 \block_reg[4][0][7]  ( .D(n2228), .CK(clk), .RN(n3741), .Q(
        \block[4][0][7] ), .QN(n607) );
  DFFRX1 \block_reg[4][0][6]  ( .D(n2229), .CK(clk), .RN(n3741), .Q(
        \block[4][0][6] ), .QN(n606) );
  DFFRX1 \block_reg[4][0][5]  ( .D(n2230), .CK(clk), .RN(n3740), .Q(
        \block[4][0][5] ), .QN(n605) );
  DFFRX1 \block_reg[4][0][4]  ( .D(n2231), .CK(clk), .RN(n3740), .Q(
        \block[4][0][4] ), .QN(n604) );
  DFFRX1 \block_reg[4][0][3]  ( .D(n2232), .CK(clk), .RN(n3740), .Q(
        \block[4][0][3] ), .QN(n603) );
  DFFRX1 \block_reg[4][0][2]  ( .D(n2233), .CK(clk), .RN(n3740), .Q(
        \block[4][0][2] ), .QN(n602) );
  DFFRX1 \block_reg[4][0][1]  ( .D(n2234), .CK(clk), .RN(n3740), .Q(
        \block[4][0][1] ), .QN(n601) );
  DFFRX1 \block_reg[4][0][0]  ( .D(n2235), .CK(clk), .RN(n3740), .Q(
        \block[4][0][0] ), .QN(n600) );
  DFFRX1 \block_reg[0][3][31]  ( .D(n2620), .CK(clk), .RN(n3735), .Q(
        \block[0][3][31] ), .QN(n1510) );
  DFFRX1 \block_reg[0][3][30]  ( .D(n2621), .CK(clk), .RN(n3735), .Q(
        \block[0][3][30] ), .QN(n1509) );
  DFFRX1 \block_reg[0][3][29]  ( .D(n2622), .CK(clk), .RN(n3734), .Q(
        \block[0][3][29] ), .QN(n1508) );
  DFFRX1 \block_reg[0][3][28]  ( .D(n2623), .CK(clk), .RN(n3734), .Q(
        \block[0][3][28] ), .QN(n1507) );
  DFFRX1 \block_reg[0][3][27]  ( .D(n2624), .CK(clk), .RN(n3734), .Q(
        \block[0][3][27] ), .QN(n1506) );
  DFFRX1 \block_reg[0][3][26]  ( .D(n2625), .CK(clk), .RN(n3734), .Q(
        \block[0][3][26] ), .QN(n1505) );
  DFFRX1 \block_reg[0][3][25]  ( .D(n2626), .CK(clk), .RN(n3734), .Q(
        \block[0][3][25] ), .QN(n1504) );
  DFFRX1 \block_reg[0][3][24]  ( .D(n2627), .CK(clk), .RN(n3734), .Q(
        \block[0][3][24] ), .QN(n1503) );
  DFFRX1 \block_reg[0][3][23]  ( .D(n2628), .CK(clk), .RN(n3734), .Q(
        \block[0][3][23] ), .QN(n1502) );
  DFFRX1 \block_reg[0][3][22]  ( .D(n2629), .CK(clk), .RN(n3734), .Q(
        \block[0][3][22] ), .QN(n1501) );
  DFFRX1 \block_reg[0][3][21]  ( .D(n2630), .CK(clk), .RN(n3734), .Q(
        \block[0][3][21] ), .QN(n1500) );
  DFFRX1 \block_reg[0][3][20]  ( .D(n2631), .CK(clk), .RN(n3734), .Q(
        \block[0][3][20] ), .QN(n1499) );
  DFFRX1 \block_reg[0][3][19]  ( .D(n2632), .CK(clk), .RN(n3734), .Q(
        \block[0][3][19] ), .QN(n1498) );
  DFFRX1 \block_reg[0][3][18]  ( .D(n2633), .CK(clk), .RN(n3734), .Q(
        \block[0][3][18] ), .QN(n1497) );
  DFFRX1 \block_reg[0][3][17]  ( .D(n2634), .CK(clk), .RN(n3733), .Q(
        \block[0][3][17] ), .QN(n1496) );
  DFFRX1 \block_reg[0][3][16]  ( .D(n2635), .CK(clk), .RN(n3733), .Q(
        \block[0][3][16] ), .QN(n1495) );
  DFFRX1 \block_reg[0][3][15]  ( .D(n2636), .CK(clk), .RN(n3733), .Q(
        \block[0][3][15] ), .QN(n1494) );
  DFFRX1 \block_reg[0][3][14]  ( .D(n2637), .CK(clk), .RN(n3733), .Q(
        \block[0][3][14] ), .QN(n1493) );
  DFFRX1 \block_reg[0][3][13]  ( .D(n2638), .CK(clk), .RN(n3733), .Q(
        \block[0][3][13] ), .QN(n1492) );
  DFFRX1 \block_reg[0][3][12]  ( .D(n2639), .CK(clk), .RN(n3733), .Q(
        \block[0][3][12] ), .QN(n1491) );
  DFFRX1 \block_reg[0][3][11]  ( .D(n2640), .CK(clk), .RN(n3733), .Q(
        \block[0][3][11] ), .QN(n1490) );
  DFFRX1 \block_reg[0][3][10]  ( .D(n2641), .CK(clk), .RN(n3733), .Q(
        \block[0][3][10] ), .QN(n1489) );
  DFFRX1 \block_reg[0][3][9]  ( .D(n2642), .CK(clk), .RN(n3733), .Q(
        \block[0][3][9] ), .QN(n1488) );
  DFFRX1 \block_reg[0][3][8]  ( .D(n2643), .CK(clk), .RN(n3733), .Q(
        \block[0][3][8] ), .QN(n1487) );
  DFFRX1 \block_reg[0][3][7]  ( .D(n2644), .CK(clk), .RN(n3733), .Q(
        \block[0][3][7] ), .QN(n1486) );
  DFFRX1 \block_reg[0][3][6]  ( .D(n2645), .CK(clk), .RN(n3733), .Q(
        \block[0][3][6] ), .QN(n1485) );
  DFFRX1 \block_reg[0][3][5]  ( .D(n2646), .CK(clk), .RN(n3732), .Q(
        \block[0][3][5] ), .QN(n1484) );
  DFFRX1 \block_reg[0][3][4]  ( .D(n2647), .CK(clk), .RN(n3732), .Q(
        \block[0][3][4] ), .QN(n1483) );
  DFFRX1 \block_reg[0][3][3]  ( .D(n2648), .CK(clk), .RN(n3732), .Q(
        \block[0][3][3] ), .QN(n1482) );
  DFFRX1 \block_reg[0][3][2]  ( .D(n2649), .CK(clk), .RN(n3732), .Q(
        \block[0][3][2] ), .QN(n1481) );
  DFFRX1 \block_reg[0][3][1]  ( .D(n2650), .CK(clk), .RN(n3732), .Q(
        \block[0][3][1] ), .QN(n1480) );
  DFFRX1 \block_reg[0][3][0]  ( .D(n2651), .CK(clk), .RN(n3732), .Q(
        \block[0][3][0] ), .QN(n1479) );
  DFFRX1 \block_reg[4][3][31]  ( .D(n2108), .CK(clk), .RN(n3724), .Q(
        \block[4][3][31] ), .QN(n727) );
  DFFRX1 \block_reg[4][3][30]  ( .D(n2109), .CK(clk), .RN(n3724), .Q(
        \block[4][3][30] ), .QN(n726) );
  DFFRX1 \block_reg[4][3][29]  ( .D(n2110), .CK(clk), .RN(n3724), .Q(
        \block[4][3][29] ), .QN(n725) );
  DFFRX1 \block_reg[4][3][28]  ( .D(n2111), .CK(clk), .RN(n3724), .Q(
        \block[4][3][28] ), .QN(n724) );
  DFFRX1 \block_reg[4][3][27]  ( .D(n2112), .CK(clk), .RN(n3724), .Q(
        \block[4][3][27] ), .QN(n723) );
  DFFRX1 \block_reg[4][3][26]  ( .D(n2113), .CK(clk), .RN(n3724), .Q(
        \block[4][3][26] ), .QN(n722) );
  DFFRX1 \block_reg[4][3][25]  ( .D(n2114), .CK(clk), .RN(n3723), .Q(
        \block[4][3][25] ), .QN(n721) );
  DFFRX1 \block_reg[4][3][24]  ( .D(n2115), .CK(clk), .RN(n3723), .Q(
        \block[4][3][24] ), .QN(n720) );
  DFFRX1 \block_reg[4][3][23]  ( .D(n2116), .CK(clk), .RN(n3723), .Q(
        \block[4][3][23] ), .QN(n719) );
  DFFRX1 \block_reg[4][3][22]  ( .D(n2117), .CK(clk), .RN(n3723), .Q(
        \block[4][3][22] ), .QN(n718) );
  DFFRX1 \block_reg[4][3][21]  ( .D(n2118), .CK(clk), .RN(n3723), .Q(
        \block[4][3][21] ), .QN(n717) );
  DFFRX1 \block_reg[4][3][20]  ( .D(n2119), .CK(clk), .RN(n3723), .Q(
        \block[4][3][20] ), .QN(n716) );
  DFFRX1 \block_reg[4][3][19]  ( .D(n2120), .CK(clk), .RN(n3723), .Q(
        \block[4][3][19] ), .QN(n715) );
  DFFRX1 \block_reg[4][3][18]  ( .D(n2121), .CK(clk), .RN(n3723), .Q(
        \block[4][3][18] ), .QN(n714) );
  DFFRX1 \block_reg[4][3][17]  ( .D(n2122), .CK(clk), .RN(n3723), .Q(
        \block[4][3][17] ), .QN(n713) );
  DFFRX1 \block_reg[4][3][16]  ( .D(n2123), .CK(clk), .RN(n3723), .Q(
        \block[4][3][16] ), .QN(n712) );
  DFFRX1 \block_reg[4][3][15]  ( .D(n2124), .CK(clk), .RN(n3723), .Q(
        \block[4][3][15] ), .QN(n711) );
  DFFRX1 \block_reg[4][3][14]  ( .D(n2125), .CK(clk), .RN(n3723), .Q(
        \block[4][3][14] ), .QN(n710) );
  DFFRX1 \block_reg[4][3][13]  ( .D(n2126), .CK(clk), .RN(n3722), .Q(
        \block[4][3][13] ), .QN(n709) );
  DFFRX1 \block_reg[4][3][12]  ( .D(n2127), .CK(clk), .RN(n3722), .Q(
        \block[4][3][12] ), .QN(n708) );
  DFFRX1 \block_reg[4][3][11]  ( .D(n2128), .CK(clk), .RN(n3722), .Q(
        \block[4][3][11] ), .QN(n707) );
  DFFRX1 \block_reg[4][3][10]  ( .D(n2129), .CK(clk), .RN(n3722), .Q(
        \block[4][3][10] ), .QN(n706) );
  DFFRX1 \block_reg[4][3][9]  ( .D(n2130), .CK(clk), .RN(n3722), .Q(
        \block[4][3][9] ), .QN(n705) );
  DFFRX1 \block_reg[4][3][8]  ( .D(n2131), .CK(clk), .RN(n3722), .Q(
        \block[4][3][8] ), .QN(n704) );
  DFFRX1 \block_reg[4][3][7]  ( .D(n2132), .CK(clk), .RN(n3722), .Q(
        \block[4][3][7] ), .QN(n703) );
  DFFRX1 \block_reg[4][3][6]  ( .D(n2133), .CK(clk), .RN(n3722), .Q(
        \block[4][3][6] ), .QN(n702) );
  DFFRX1 \block_reg[4][3][5]  ( .D(n2134), .CK(clk), .RN(n3722), .Q(
        \block[4][3][5] ), .QN(n701) );
  DFFRX1 \block_reg[4][3][4]  ( .D(n2135), .CK(clk), .RN(n3722), .Q(
        \block[4][3][4] ), .QN(n700) );
  DFFRX1 \block_reg[4][3][3]  ( .D(n2136), .CK(clk), .RN(n3722), .Q(
        \block[4][3][3] ), .QN(n699) );
  DFFRX1 \block_reg[4][3][2]  ( .D(n2137), .CK(clk), .RN(n3722), .Q(
        \block[4][3][2] ), .QN(n698) );
  DFFRX1 \block_reg[4][3][1]  ( .D(n2138), .CK(clk), .RN(n3721), .Q(
        \block[4][3][1] ), .QN(n697) );
  DFFRX1 \block_reg[4][3][0]  ( .D(n2139), .CK(clk), .RN(n3721), .Q(
        \block[4][3][0] ), .QN(n696) );
  DFFRX1 \block_reg[0][2][31]  ( .D(n2652), .CK(clk), .RN(n3713), .Q(
        \block[0][2][31] ), .QN(n1478) );
  DFFRX1 \block_reg[0][2][30]  ( .D(n2653), .CK(clk), .RN(n3713), .Q(
        \block[0][2][30] ), .QN(n1477) );
  DFFRX1 \block_reg[0][2][29]  ( .D(n2654), .CK(clk), .RN(n3713), .Q(
        \block[0][2][29] ), .QN(n1476) );
  DFFRX1 \block_reg[0][2][28]  ( .D(n2655), .CK(clk), .RN(n3713), .Q(
        \block[0][2][28] ), .QN(n1475) );
  DFFRX1 \block_reg[0][2][27]  ( .D(n2656), .CK(clk), .RN(n3713), .Q(
        \block[0][2][27] ), .QN(n1474) );
  DFFRX1 \block_reg[0][2][26]  ( .D(n2657), .CK(clk), .RN(n3713), .Q(
        \block[0][2][26] ), .QN(n1473) );
  DFFRX1 \block_reg[0][2][25]  ( .D(n2658), .CK(clk), .RN(n3713), .Q(
        \block[0][2][25] ), .QN(n1472) );
  DFFRX1 \block_reg[0][2][24]  ( .D(n2659), .CK(clk), .RN(n3713), .Q(
        \block[0][2][24] ), .QN(n1471) );
  DFFRX1 \block_reg[0][2][23]  ( .D(n2660), .CK(clk), .RN(n3713), .Q(
        \block[0][2][23] ), .QN(n1470) );
  DFFRX1 \block_reg[0][2][22]  ( .D(n2661), .CK(clk), .RN(n3713), .Q(
        \block[0][2][22] ), .QN(n1469) );
  DFFRX1 \block_reg[0][2][21]  ( .D(n2662), .CK(clk), .RN(n3712), .Q(
        \block[0][2][21] ), .QN(n1468) );
  DFFRX1 \block_reg[0][2][20]  ( .D(n2663), .CK(clk), .RN(n3712), .Q(
        \block[0][2][20] ), .QN(n1467) );
  DFFRX1 \block_reg[0][2][19]  ( .D(n2664), .CK(clk), .RN(n3712), .Q(
        \block[0][2][19] ), .QN(n1466) );
  DFFRX1 \block_reg[0][2][18]  ( .D(n2665), .CK(clk), .RN(n3712), .Q(
        \block[0][2][18] ), .QN(n1465) );
  DFFRX1 \block_reg[0][2][17]  ( .D(n2666), .CK(clk), .RN(n3712), .Q(
        \block[0][2][17] ), .QN(n1464) );
  DFFRX1 \block_reg[0][2][16]  ( .D(n2667), .CK(clk), .RN(n3712), .Q(
        \block[0][2][16] ), .QN(n1463) );
  DFFRX1 \block_reg[0][2][15]  ( .D(n2668), .CK(clk), .RN(n3712), .Q(
        \block[0][2][15] ), .QN(n1462) );
  DFFRX1 \block_reg[0][2][14]  ( .D(n2669), .CK(clk), .RN(n3712), .Q(
        \block[0][2][14] ), .QN(n1461) );
  DFFRX1 \block_reg[0][2][13]  ( .D(n2670), .CK(clk), .RN(n3712), .Q(
        \block[0][2][13] ), .QN(n1460) );
  DFFRX1 \block_reg[0][2][12]  ( .D(n2671), .CK(clk), .RN(n3712), .Q(
        \block[0][2][12] ), .QN(n1459) );
  DFFRX1 \block_reg[0][2][11]  ( .D(n2672), .CK(clk), .RN(n3712), .Q(
        \block[0][2][11] ), .QN(n1458) );
  DFFRX1 \block_reg[0][2][10]  ( .D(n2673), .CK(clk), .RN(n3712), .Q(
        \block[0][2][10] ), .QN(n1457) );
  DFFRX1 \block_reg[0][2][9]  ( .D(n2674), .CK(clk), .RN(n3711), .Q(
        \block[0][2][9] ), .QN(n1456) );
  DFFRX1 \block_reg[0][2][8]  ( .D(n2675), .CK(clk), .RN(n3711), .Q(
        \block[0][2][8] ), .QN(n1455) );
  DFFRX1 \block_reg[0][2][7]  ( .D(n2676), .CK(clk), .RN(n3711), .Q(
        \block[0][2][7] ), .QN(n1454) );
  DFFRX1 \block_reg[0][2][6]  ( .D(n2677), .CK(clk), .RN(n3711), .Q(
        \block[0][2][6] ), .QN(n1453) );
  DFFRX1 \block_reg[0][2][5]  ( .D(n2678), .CK(clk), .RN(n3711), .Q(
        \block[0][2][5] ), .QN(n1452) );
  DFFRX1 \block_reg[0][2][4]  ( .D(n2679), .CK(clk), .RN(n3711), .Q(
        \block[0][2][4] ), .QN(n1451) );
  DFFRX1 \block_reg[0][2][3]  ( .D(n2680), .CK(clk), .RN(n3711), .Q(
        \block[0][2][3] ), .QN(n1450) );
  DFFRX1 \block_reg[0][2][2]  ( .D(n2681), .CK(clk), .RN(n3711), .Q(
        \block[0][2][2] ), .QN(n1449) );
  DFFRX1 \block_reg[0][2][1]  ( .D(n2682), .CK(clk), .RN(n3711), .Q(
        \block[0][2][1] ), .QN(n1448) );
  DFFRX1 \block_reg[0][2][0]  ( .D(n2683), .CK(clk), .RN(n3711), .Q(
        \block[0][2][0] ), .QN(n1447) );
  DFFRX1 \block_reg[4][2][31]  ( .D(n2140), .CK(clk), .RN(n3703), .Q(
        \block[4][2][31] ), .QN(n695) );
  DFFRX1 \block_reg[4][2][30]  ( .D(n2141), .CK(clk), .RN(n3703), .Q(
        \block[4][2][30] ), .QN(n694) );
  DFFRX1 \block_reg[4][2][29]  ( .D(n2142), .CK(clk), .RN(n3702), .Q(
        \block[4][2][29] ), .QN(n693) );
  DFFRX1 \block_reg[4][2][28]  ( .D(n2143), .CK(clk), .RN(n3702), .Q(
        \block[4][2][28] ), .QN(n692) );
  DFFRX1 \block_reg[4][2][27]  ( .D(n2144), .CK(clk), .RN(n3702), .Q(
        \block[4][2][27] ), .QN(n691) );
  DFFRX1 \block_reg[4][2][26]  ( .D(n2145), .CK(clk), .RN(n3702), .Q(
        \block[4][2][26] ), .QN(n690) );
  DFFRX1 \block_reg[4][2][25]  ( .D(n2146), .CK(clk), .RN(n3702), .Q(
        \block[4][2][25] ), .QN(n689) );
  DFFRX1 \block_reg[4][2][24]  ( .D(n2147), .CK(clk), .RN(n3702), .Q(
        \block[4][2][24] ), .QN(n688) );
  DFFRX1 \block_reg[4][2][23]  ( .D(n2148), .CK(clk), .RN(n3702), .Q(
        \block[4][2][23] ), .QN(n687) );
  DFFRX1 \block_reg[4][2][22]  ( .D(n2149), .CK(clk), .RN(n3702), .Q(
        \block[4][2][22] ), .QN(n686) );
  DFFRX1 \block_reg[4][2][21]  ( .D(n2150), .CK(clk), .RN(n3702), .Q(
        \block[4][2][21] ), .QN(n685) );
  DFFRX1 \block_reg[4][2][20]  ( .D(n2151), .CK(clk), .RN(n3702), .Q(
        \block[4][2][20] ), .QN(n684) );
  DFFRX1 \block_reg[4][2][19]  ( .D(n2152), .CK(clk), .RN(n3702), .Q(
        \block[4][2][19] ), .QN(n683) );
  DFFRX1 \block_reg[4][2][18]  ( .D(n2153), .CK(clk), .RN(n3702), .Q(
        \block[4][2][18] ), .QN(n682) );
  DFFRX1 \block_reg[4][2][17]  ( .D(n2154), .CK(clk), .RN(n3701), .Q(
        \block[4][2][17] ), .QN(n681) );
  DFFRX1 \block_reg[4][2][16]  ( .D(n2155), .CK(clk), .RN(n3701), .Q(
        \block[4][2][16] ), .QN(n680) );
  DFFRX1 \block_reg[4][2][15]  ( .D(n2156), .CK(clk), .RN(n3701), .Q(
        \block[4][2][15] ), .QN(n679) );
  DFFRX1 \block_reg[4][2][14]  ( .D(n2157), .CK(clk), .RN(n3701), .Q(
        \block[4][2][14] ), .QN(n678) );
  DFFRX1 \block_reg[4][2][13]  ( .D(n2158), .CK(clk), .RN(n3701), .Q(
        \block[4][2][13] ), .QN(n677) );
  DFFRX1 \block_reg[4][2][12]  ( .D(n2159), .CK(clk), .RN(n3701), .Q(
        \block[4][2][12] ), .QN(n676) );
  DFFRX1 \block_reg[4][2][11]  ( .D(n2160), .CK(clk), .RN(n3701), .Q(
        \block[4][2][11] ), .QN(n675) );
  DFFRX1 \block_reg[4][2][10]  ( .D(n2161), .CK(clk), .RN(n3701), .Q(
        \block[4][2][10] ), .QN(n674) );
  DFFRX1 \block_reg[4][2][9]  ( .D(n2162), .CK(clk), .RN(n3701), .Q(
        \block[4][2][9] ), .QN(n673) );
  DFFRX1 \block_reg[4][2][8]  ( .D(n2163), .CK(clk), .RN(n3701), .Q(
        \block[4][2][8] ), .QN(n672) );
  DFFRX1 \block_reg[4][2][7]  ( .D(n2164), .CK(clk), .RN(n3701), .Q(
        \block[4][2][7] ), .QN(n671) );
  DFFRX1 \block_reg[4][2][6]  ( .D(n2165), .CK(clk), .RN(n3701), .Q(
        \block[4][2][6] ), .QN(n670) );
  DFFRX1 \block_reg[4][2][5]  ( .D(n2166), .CK(clk), .RN(n3700), .Q(
        \block[4][2][5] ), .QN(n669) );
  DFFRX1 \block_reg[4][2][4]  ( .D(n2167), .CK(clk), .RN(n3700), .Q(
        \block[4][2][4] ), .QN(n668) );
  DFFRX1 \block_reg[4][2][3]  ( .D(n2168), .CK(clk), .RN(n3700), .Q(
        \block[4][2][3] ), .QN(n667) );
  DFFRX1 \block_reg[4][2][2]  ( .D(n2169), .CK(clk), .RN(n3700), .Q(
        \block[4][2][2] ), .QN(n666) );
  DFFRX1 \block_reg[4][2][1]  ( .D(n2170), .CK(clk), .RN(n3700), .Q(
        \block[4][2][1] ), .QN(n665) );
  DFFRX1 \block_reg[4][2][0]  ( .D(n2171), .CK(clk), .RN(n3700), .Q(
        \block[4][2][0] ), .QN(n664) );
  DFFRX1 \block_reg[0][1][31]  ( .D(n2684), .CK(clk), .RN(n3692), .Q(
        \block[0][1][31] ), .QN(n1446) );
  DFFRX1 \block_reg[0][1][30]  ( .D(n2685), .CK(clk), .RN(n3692), .Q(
        \block[0][1][30] ), .QN(n1445) );
  DFFRX1 \block_reg[0][1][29]  ( .D(n2686), .CK(clk), .RN(n3692), .Q(
        \block[0][1][29] ), .QN(n1444) );
  DFFRX1 \block_reg[0][1][28]  ( .D(n2687), .CK(clk), .RN(n3692), .Q(
        \block[0][1][28] ), .QN(n1443) );
  DFFRX1 \block_reg[0][1][27]  ( .D(n2688), .CK(clk), .RN(n3692), .Q(
        \block[0][1][27] ), .QN(n1442) );
  DFFRX1 \block_reg[0][1][26]  ( .D(n2689), .CK(clk), .RN(n3692), .Q(
        \block[0][1][26] ), .QN(n1441) );
  DFFRX1 \block_reg[0][1][25]  ( .D(n2690), .CK(clk), .RN(n3691), .Q(
        \block[0][1][25] ), .QN(n1440) );
  DFFRX1 \block_reg[0][1][24]  ( .D(n2691), .CK(clk), .RN(n3691), .Q(
        \block[0][1][24] ), .QN(n1439) );
  DFFRX1 \block_reg[0][1][23]  ( .D(n2692), .CK(clk), .RN(n3691), .Q(
        \block[0][1][23] ), .QN(n1438) );
  DFFRX1 \block_reg[0][1][22]  ( .D(n2693), .CK(clk), .RN(n3691), .Q(
        \block[0][1][22] ), .QN(n1437) );
  DFFRX1 \block_reg[0][1][21]  ( .D(n2694), .CK(clk), .RN(n3691), .Q(
        \block[0][1][21] ), .QN(n1436) );
  DFFRX1 \block_reg[0][1][20]  ( .D(n2695), .CK(clk), .RN(n3691), .Q(
        \block[0][1][20] ), .QN(n1435) );
  DFFRX1 \block_reg[0][1][19]  ( .D(n2696), .CK(clk), .RN(n3691), .Q(
        \block[0][1][19] ), .QN(n1434) );
  DFFRX1 \block_reg[0][1][18]  ( .D(n2697), .CK(clk), .RN(n3691), .Q(
        \block[0][1][18] ), .QN(n1433) );
  DFFRX1 \block_reg[0][1][17]  ( .D(n2698), .CK(clk), .RN(n3691), .Q(
        \block[0][1][17] ), .QN(n1432) );
  DFFRX1 \block_reg[0][1][16]  ( .D(n2699), .CK(clk), .RN(n3691), .Q(
        \block[0][1][16] ), .QN(n1431) );
  DFFRX1 \block_reg[0][1][15]  ( .D(n2700), .CK(clk), .RN(n3691), .Q(
        \block[0][1][15] ), .QN(n1430) );
  DFFRX1 \block_reg[0][1][14]  ( .D(n2701), .CK(clk), .RN(n3691), .Q(
        \block[0][1][14] ), .QN(n1429) );
  DFFRX1 \block_reg[0][1][13]  ( .D(n2702), .CK(clk), .RN(n3690), .Q(
        \block[0][1][13] ), .QN(n1428) );
  DFFRX1 \block_reg[0][1][12]  ( .D(n2703), .CK(clk), .RN(n3690), .Q(
        \block[0][1][12] ), .QN(n1427) );
  DFFRX1 \block_reg[0][1][11]  ( .D(n2704), .CK(clk), .RN(n3690), .Q(
        \block[0][1][11] ), .QN(n1426) );
  DFFRX1 \block_reg[0][1][10]  ( .D(n2705), .CK(clk), .RN(n3690), .Q(
        \block[0][1][10] ), .QN(n1425) );
  DFFRX1 \block_reg[0][1][9]  ( .D(n2706), .CK(clk), .RN(n3690), .Q(
        \block[0][1][9] ), .QN(n1424) );
  DFFRX1 \block_reg[0][1][8]  ( .D(n2707), .CK(clk), .RN(n3690), .Q(
        \block[0][1][8] ), .QN(n1423) );
  DFFRX1 \block_reg[0][1][7]  ( .D(n2708), .CK(clk), .RN(n3690), .Q(
        \block[0][1][7] ), .QN(n1422) );
  DFFRX1 \block_reg[0][1][6]  ( .D(n2709), .CK(clk), .RN(n3690), .Q(
        \block[0][1][6] ), .QN(n1421) );
  DFFRX1 \block_reg[0][1][5]  ( .D(n2710), .CK(clk), .RN(n3690), .Q(
        \block[0][1][5] ), .QN(n1420) );
  DFFRX1 \block_reg[0][1][4]  ( .D(n2711), .CK(clk), .RN(n3690), .Q(
        \block[0][1][4] ), .QN(n1419) );
  DFFRX1 \block_reg[0][1][3]  ( .D(n2712), .CK(clk), .RN(n3690), .Q(
        \block[0][1][3] ), .QN(n1418) );
  DFFRX1 \block_reg[0][1][2]  ( .D(n2713), .CK(clk), .RN(n3690), .Q(
        \block[0][1][2] ), .QN(n1417) );
  DFFRX1 \block_reg[0][1][1]  ( .D(n2714), .CK(clk), .RN(n3689), .Q(
        \block[0][1][1] ), .QN(n1416) );
  DFFRX1 \block_reg[0][1][0]  ( .D(n2715), .CK(clk), .RN(n3689), .Q(
        \block[0][1][0] ), .QN(n1415) );
  DFFRX1 \block_reg[4][1][31]  ( .D(n2172), .CK(clk), .RN(n3681), .Q(
        \block[4][1][31] ), .QN(n663) );
  DFFRX1 \block_reg[4][1][30]  ( .D(n2173), .CK(clk), .RN(n3681), .Q(
        \block[4][1][30] ), .QN(n662) );
  DFFRX1 \block_reg[4][1][29]  ( .D(n2174), .CK(clk), .RN(n3681), .Q(
        \block[4][1][29] ), .QN(n661) );
  DFFRX1 \block_reg[4][1][28]  ( .D(n2175), .CK(clk), .RN(n3681), .Q(
        \block[4][1][28] ), .QN(n660) );
  DFFRX1 \block_reg[4][1][27]  ( .D(n2176), .CK(clk), .RN(n3681), .Q(
        \block[4][1][27] ), .QN(n659) );
  DFFRX1 \block_reg[4][1][26]  ( .D(n2177), .CK(clk), .RN(n3681), .Q(
        \block[4][1][26] ), .QN(n658) );
  DFFRX1 \block_reg[4][1][25]  ( .D(n2178), .CK(clk), .RN(n3681), .Q(
        \block[4][1][25] ), .QN(n657) );
  DFFRX1 \block_reg[4][1][24]  ( .D(n2179), .CK(clk), .RN(n3681), .Q(
        \block[4][1][24] ), .QN(n656) );
  DFFRX1 \block_reg[4][1][23]  ( .D(n2180), .CK(clk), .RN(n3681), .Q(
        \block[4][1][23] ), .QN(n655) );
  DFFRX1 \block_reg[4][1][22]  ( .D(n2181), .CK(clk), .RN(n3681), .Q(
        \block[4][1][22] ), .QN(n654) );
  DFFRX1 \block_reg[4][1][21]  ( .D(n2182), .CK(clk), .RN(n3680), .Q(
        \block[4][1][21] ), .QN(n653) );
  DFFRX1 \block_reg[4][1][20]  ( .D(n2183), .CK(clk), .RN(n3680), .Q(
        \block[4][1][20] ), .QN(n652) );
  DFFRX1 \block_reg[4][1][19]  ( .D(n2184), .CK(clk), .RN(n3680), .Q(
        \block[4][1][19] ), .QN(n651) );
  DFFRX1 \block_reg[4][1][18]  ( .D(n2185), .CK(clk), .RN(n3680), .Q(
        \block[4][1][18] ), .QN(n650) );
  DFFRX1 \block_reg[4][1][17]  ( .D(n2186), .CK(clk), .RN(n3680), .Q(
        \block[4][1][17] ), .QN(n649) );
  DFFRX1 \block_reg[4][1][16]  ( .D(n2187), .CK(clk), .RN(n3680), .Q(
        \block[4][1][16] ), .QN(n648) );
  DFFRX1 \block_reg[4][1][15]  ( .D(n2188), .CK(clk), .RN(n3680), .Q(
        \block[4][1][15] ), .QN(n647) );
  DFFRX1 \block_reg[4][1][14]  ( .D(n2189), .CK(clk), .RN(n3680), .Q(
        \block[4][1][14] ), .QN(n646) );
  DFFRX1 \block_reg[4][1][13]  ( .D(n2190), .CK(clk), .RN(n3680), .Q(
        \block[4][1][13] ), .QN(n645) );
  DFFRX1 \block_reg[4][1][12]  ( .D(n2191), .CK(clk), .RN(n3680), .Q(
        \block[4][1][12] ), .QN(n644) );
  DFFRX1 \block_reg[4][1][11]  ( .D(n2192), .CK(clk), .RN(n3680), .Q(
        \block[4][1][11] ), .QN(n643) );
  DFFRX1 \block_reg[4][1][10]  ( .D(n2193), .CK(clk), .RN(n3680), .Q(
        \block[4][1][10] ), .QN(n642) );
  DFFRX1 \block_reg[4][1][9]  ( .D(n2194), .CK(clk), .RN(n3679), .Q(
        \block[4][1][9] ), .QN(n641) );
  DFFRX1 \block_reg[4][1][8]  ( .D(n2195), .CK(clk), .RN(n3679), .Q(
        \block[4][1][8] ), .QN(n640) );
  DFFRX1 \block_reg[4][1][7]  ( .D(n2196), .CK(clk), .RN(n3679), .Q(
        \block[4][1][7] ), .QN(n639) );
  DFFRX1 \block_reg[4][1][6]  ( .D(n2197), .CK(clk), .RN(n3679), .Q(
        \block[4][1][6] ), .QN(n638) );
  DFFRX1 \block_reg[4][1][5]  ( .D(n2198), .CK(clk), .RN(n3679), .Q(
        \block[4][1][5] ), .QN(n637) );
  DFFRX1 \block_reg[4][1][4]  ( .D(n2199), .CK(clk), .RN(n3679), .Q(
        \block[4][1][4] ), .QN(n636) );
  DFFRX1 \block_reg[4][1][3]  ( .D(n2200), .CK(clk), .RN(n3679), .Q(
        \block[4][1][3] ), .QN(n635) );
  DFFRX1 \block_reg[4][1][2]  ( .D(n2201), .CK(clk), .RN(n3679), .Q(
        \block[4][1][2] ), .QN(n634) );
  DFFRX1 \block_reg[4][1][1]  ( .D(n2202), .CK(clk), .RN(n3679), .Q(
        \block[4][1][1] ), .QN(n633) );
  DFFRX1 \block_reg[4][1][0]  ( .D(n2203), .CK(clk), .RN(n3679), .Q(
        \block[4][1][0] ), .QN(n632) );
  DFFRX1 \dirty_reg[6]  ( .D(n1717), .CK(clk), .RN(n3759), .Q(dirty[6]), .QN(
        n1118) );
  DFFRX1 \dirty_reg[2]  ( .D(n1721), .CK(clk), .RN(n3759), .Q(dirty[2]), .QN(
        n1114) );
  DFFRX1 \valid_reg[7]  ( .D(n1711), .CK(clk), .RN(n3780), .Q(valid[7]), .QN(
        n1696) );
  DFFRX1 \tag_reg[7][24]  ( .D(n2970), .CK(clk), .RN(n3780), .Q(\tag[7][24] ), 
        .QN(n1321) );
  DFFRX1 \tag_reg[7][23]  ( .D(n2971), .CK(clk), .RN(n3780), .Q(\tag[7][23] ), 
        .QN(n1320) );
  DFFRX1 \tag_reg[7][22]  ( .D(n2972), .CK(clk), .RN(n3780), .Q(\tag[7][22] ), 
        .QN(n1319) );
  DFFRX1 \tag_reg[7][21]  ( .D(n2973), .CK(clk), .RN(n3780), .Q(\tag[7][21] ), 
        .QN(n1318) );
  DFFRX1 \tag_reg[7][20]  ( .D(n2974), .CK(clk), .RN(n3780), .QN(n1317) );
  DFFRX1 \tag_reg[7][19]  ( .D(n2975), .CK(clk), .RN(n3780), .QN(n1316) );
  DFFRX1 \tag_reg[7][18]  ( .D(n2976), .CK(clk), .RN(n3780), .Q(\tag[7][18] ), 
        .QN(n1315) );
  DFFRX1 \tag_reg[7][17]  ( .D(n2977), .CK(clk), .RN(n3780), .QN(n1314) );
  DFFRX1 \tag_reg[7][16]  ( .D(n2978), .CK(clk), .RN(n3780), .Q(\tag[7][16] ), 
        .QN(n1313) );
  DFFRX1 \tag_reg[7][15]  ( .D(n2979), .CK(clk), .RN(n3780), .Q(\tag[7][15] ), 
        .QN(n1312) );
  DFFRX1 \tag_reg[7][14]  ( .D(n2980), .CK(clk), .RN(n3780), .Q(\tag[7][14] ), 
        .QN(n1311) );
  DFFRX1 \tag_reg[7][13]  ( .D(n2981), .CK(clk), .RN(n3779), .Q(\tag[7][13] ), 
        .QN(n1310) );
  DFFRX1 \tag_reg[7][12]  ( .D(n2982), .CK(clk), .RN(n3779), .Q(\tag[7][12] ), 
        .QN(n1309) );
  DFFRX1 \tag_reg[7][11]  ( .D(n2983), .CK(clk), .RN(n3779), .Q(\tag[7][11] ), 
        .QN(n1308) );
  DFFRX1 \tag_reg[7][10]  ( .D(n2984), .CK(clk), .RN(n3779), .Q(\tag[7][10] ), 
        .QN(n1307) );
  DFFRX1 \tag_reg[7][9]  ( .D(n2985), .CK(clk), .RN(n3779), .Q(\tag[7][9] ), 
        .QN(n1306) );
  DFFRX1 \tag_reg[7][8]  ( .D(n2986), .CK(clk), .RN(n3779), .Q(\tag[7][8] ), 
        .QN(n1305) );
  DFFRX1 \tag_reg[7][7]  ( .D(n2987), .CK(clk), .RN(n3779), .QN(n1304) );
  DFFRX1 \tag_reg[7][6]  ( .D(n2988), .CK(clk), .RN(n3779), .QN(n1303) );
  DFFRX1 \tag_reg[7][5]  ( .D(n2989), .CK(clk), .RN(n3779), .QN(n1302) );
  DFFRX1 \tag_reg[7][4]  ( .D(n2990), .CK(clk), .RN(n3779), .QN(n1301) );
  DFFRX1 \tag_reg[7][3]  ( .D(n2991), .CK(clk), .RN(n3779), .Q(\tag[7][3] ), 
        .QN(n1300) );
  DFFRX1 \tag_reg[7][2]  ( .D(n2992), .CK(clk), .RN(n3779), .QN(n1299) );
  DFFRX1 \tag_reg[7][1]  ( .D(n2993), .CK(clk), .RN(n3778), .Q(\tag[7][1] ), 
        .QN(n1298) );
  DFFRX1 \tag_reg[7][0]  ( .D(n2994), .CK(clk), .RN(n3778), .Q(\tag[7][0] ), 
        .QN(n1297) );
  DFFRX1 \valid_reg[3]  ( .D(n1707), .CK(clk), .RN(n3772), .Q(valid[3]), .QN(
        n1700) );
  DFFRX1 \tag_reg[3][24]  ( .D(n3070), .CK(clk), .RN(n3772), .Q(\tag[3][24] ), 
        .QN(n1221) );
  DFFRX1 \tag_reg[3][23]  ( .D(n3071), .CK(clk), .RN(n3772), .Q(\tag[3][23] ), 
        .QN(n1220) );
  DFFRX1 \tag_reg[3][22]  ( .D(n3072), .CK(clk), .RN(n3772), .Q(\tag[3][22] ), 
        .QN(n1219) );
  DFFRX1 \tag_reg[3][21]  ( .D(n3073), .CK(clk), .RN(n3771), .Q(\tag[3][21] ), 
        .QN(n1218) );
  DFFRX1 \tag_reg[3][20]  ( .D(n3074), .CK(clk), .RN(n3771), .QN(n1217) );
  DFFRX1 \tag_reg[3][19]  ( .D(n3075), .CK(clk), .RN(n3771), .QN(n1216) );
  DFFRX1 \tag_reg[3][18]  ( .D(n3076), .CK(clk), .RN(n3771), .Q(\tag[3][18] ), 
        .QN(n1215) );
  DFFRX1 \tag_reg[3][17]  ( .D(n3077), .CK(clk), .RN(n3771), .QN(n1214) );
  DFFRX1 \tag_reg[3][16]  ( .D(n3078), .CK(clk), .RN(n3771), .Q(\tag[3][16] ), 
        .QN(n1213) );
  DFFRX1 \tag_reg[3][15]  ( .D(n3079), .CK(clk), .RN(n3771), .Q(\tag[3][15] ), 
        .QN(n1212) );
  DFFRX1 \tag_reg[3][14]  ( .D(n3080), .CK(clk), .RN(n3771), .Q(\tag[3][14] ), 
        .QN(n1211) );
  DFFRX1 \tag_reg[3][13]  ( .D(n3081), .CK(clk), .RN(n3771), .Q(\tag[3][13] ), 
        .QN(n1210) );
  DFFRX1 \tag_reg[3][12]  ( .D(n3082), .CK(clk), .RN(n3771), .Q(\tag[3][12] ), 
        .QN(n1209) );
  DFFRX1 \tag_reg[3][11]  ( .D(n3083), .CK(clk), .RN(n3771), .Q(\tag[3][11] ), 
        .QN(n1208) );
  DFFRX1 \tag_reg[3][10]  ( .D(n3084), .CK(clk), .RN(n3771), .Q(\tag[3][10] ), 
        .QN(n1207) );
  DFFRX1 \tag_reg[3][9]  ( .D(n3085), .CK(clk), .RN(n3770), .Q(\tag[3][9] ), 
        .QN(n1206) );
  DFFRX1 \tag_reg[3][8]  ( .D(n3086), .CK(clk), .RN(n3770), .Q(\tag[3][8] ), 
        .QN(n1205) );
  DFFRX1 \tag_reg[3][7]  ( .D(n3087), .CK(clk), .RN(n3770), .QN(n1204) );
  DFFRX1 \tag_reg[3][6]  ( .D(n3088), .CK(clk), .RN(n3770), .QN(n1203) );
  DFFRX1 \tag_reg[3][5]  ( .D(n3089), .CK(clk), .RN(n3770), .QN(n1202) );
  DFFRX1 \tag_reg[3][4]  ( .D(n3090), .CK(clk), .RN(n3770), .QN(n1201) );
  DFFRX1 \tag_reg[3][3]  ( .D(n3091), .CK(clk), .RN(n3770), .Q(\tag[3][3] ), 
        .QN(n1200) );
  DFFRX1 \tag_reg[3][2]  ( .D(n3092), .CK(clk), .RN(n3770), .QN(n1199) );
  DFFRX1 \tag_reg[3][1]  ( .D(n3093), .CK(clk), .RN(n3770), .Q(\tag[3][1] ), 
        .QN(n1198) );
  DFFRX1 \tag_reg[3][0]  ( .D(n3094), .CK(clk), .RN(n3770), .Q(\tag[3][0] ), 
        .QN(n1197) );
  DFFRX1 \valid_reg[5]  ( .D(n1709), .CK(clk), .RN(n3776), .Q(valid[5]), .QN(
        n1698) );
  DFFRX1 \tag_reg[5][24]  ( .D(n3020), .CK(clk), .RN(n3776), .Q(\tag[5][24] ), 
        .QN(n1271) );
  DFFRX1 \tag_reg[5][23]  ( .D(n3021), .CK(clk), .RN(n3776), .Q(\tag[5][23] ), 
        .QN(n1270) );
  DFFRX1 \tag_reg[5][22]  ( .D(n3022), .CK(clk), .RN(n3776), .Q(\tag[5][22] ), 
        .QN(n1269) );
  DFFRX1 \tag_reg[5][21]  ( .D(n3023), .CK(clk), .RN(n3776), .Q(\tag[5][21] ), 
        .QN(n1268) );
  DFFRX1 \tag_reg[5][20]  ( .D(n3024), .CK(clk), .RN(n3776), .QN(n1267) );
  DFFRX1 \tag_reg[5][19]  ( .D(n3025), .CK(clk), .RN(n3776), .QN(n1266) );
  DFFRX1 \tag_reg[5][18]  ( .D(n3026), .CK(clk), .RN(n3776), .Q(\tag[5][18] ), 
        .QN(n1265) );
  DFFRX1 \tag_reg[5][17]  ( .D(n3027), .CK(clk), .RN(n3775), .QN(n1264) );
  DFFRX1 \tag_reg[5][16]  ( .D(n3028), .CK(clk), .RN(n3775), .Q(\tag[5][16] ), 
        .QN(n1263) );
  DFFRX1 \tag_reg[5][15]  ( .D(n3029), .CK(clk), .RN(n3775), .Q(\tag[5][15] ), 
        .QN(n1262) );
  DFFRX1 \tag_reg[5][14]  ( .D(n3030), .CK(clk), .RN(n3775), .Q(\tag[5][14] ), 
        .QN(n1261) );
  DFFRX1 \tag_reg[5][13]  ( .D(n3031), .CK(clk), .RN(n3775), .Q(\tag[5][13] ), 
        .QN(n1260) );
  DFFRX1 \tag_reg[5][12]  ( .D(n3032), .CK(clk), .RN(n3775), .Q(\tag[5][12] ), 
        .QN(n1259) );
  DFFRX1 \tag_reg[5][11]  ( .D(n3033), .CK(clk), .RN(n3775), .Q(\tag[5][11] ), 
        .QN(n1258) );
  DFFRX1 \tag_reg[5][10]  ( .D(n3034), .CK(clk), .RN(n3775), .Q(\tag[5][10] ), 
        .QN(n1257) );
  DFFRX1 \tag_reg[5][9]  ( .D(n3035), .CK(clk), .RN(n3775), .Q(\tag[5][9] ), 
        .QN(n1256) );
  DFFRX1 \tag_reg[5][8]  ( .D(n3036), .CK(clk), .RN(n3775), .Q(\tag[5][8] ), 
        .QN(n1255) );
  DFFRX1 \tag_reg[5][7]  ( .D(n3037), .CK(clk), .RN(n3775), .QN(n1254) );
  DFFRX1 \tag_reg[5][6]  ( .D(n3038), .CK(clk), .RN(n3775), .QN(n1253) );
  DFFRX1 \tag_reg[5][5]  ( .D(n3039), .CK(clk), .RN(n3774), .QN(n1252) );
  DFFRX1 \tag_reg[5][4]  ( .D(n3040), .CK(clk), .RN(n3774), .QN(n1251) );
  DFFRX1 \tag_reg[5][3]  ( .D(n3041), .CK(clk), .RN(n3774), .Q(\tag[5][3] ), 
        .QN(n1250) );
  DFFRX1 \tag_reg[5][2]  ( .D(n3042), .CK(clk), .RN(n3774), .QN(n1249) );
  DFFRX1 \tag_reg[5][1]  ( .D(n3043), .CK(clk), .RN(n3774), .Q(\tag[5][1] ), 
        .QN(n1248) );
  DFFRX1 \tag_reg[5][0]  ( .D(n3044), .CK(clk), .RN(n3774), .Q(\tag[5][0] ), 
        .QN(n1247) );
  DFFRX1 \valid_reg[1]  ( .D(n1705), .CK(clk), .RN(n3767), .Q(valid[1]), .QN(
        n1702) );
  DFFRX1 \tag_reg[1][24]  ( .D(n3120), .CK(clk), .RN(n3767), .Q(\tag[1][24] ), 
        .QN(n1171) );
  DFFRX1 \tag_reg[1][23]  ( .D(n3121), .CK(clk), .RN(n3767), .Q(\tag[1][23] ), 
        .QN(n1170) );
  DFFRX1 \tag_reg[1][22]  ( .D(n3122), .CK(clk), .RN(n3767), .Q(\tag[1][22] ), 
        .QN(n1169) );
  DFFRX1 \tag_reg[1][21]  ( .D(n3123), .CK(clk), .RN(n3767), .Q(\tag[1][21] ), 
        .QN(n1168) );
  DFFRX1 \tag_reg[1][20]  ( .D(n3124), .CK(clk), .RN(n3767), .QN(n1167) );
  DFFRX1 \tag_reg[1][19]  ( .D(n3125), .CK(clk), .RN(n3767), .QN(n1166) );
  DFFRX1 \tag_reg[1][18]  ( .D(n3126), .CK(clk), .RN(n3767), .Q(\tag[1][18] ), 
        .QN(n1165) );
  DFFRX1 \tag_reg[1][17]  ( .D(n3127), .CK(clk), .RN(n3767), .QN(n1164) );
  DFFRX1 \tag_reg[1][16]  ( .D(n3128), .CK(clk), .RN(n3767), .Q(\tag[1][16] ), 
        .QN(n1163) );
  DFFRX1 \tag_reg[1][15]  ( .D(n3129), .CK(clk), .RN(n3767), .Q(\tag[1][15] ), 
        .QN(n1162) );
  DFFRX1 \tag_reg[1][14]  ( .D(n3130), .CK(clk), .RN(n3767), .Q(\tag[1][14] ), 
        .QN(n1161) );
  DFFRX1 \tag_reg[1][13]  ( .D(n3131), .CK(clk), .RN(n3766), .Q(\tag[1][13] ), 
        .QN(n1160) );
  DFFRX1 \tag_reg[1][12]  ( .D(n3132), .CK(clk), .RN(n3766), .Q(\tag[1][12] ), 
        .QN(n1159) );
  DFFRX1 \tag_reg[1][11]  ( .D(n3133), .CK(clk), .RN(n3766), .Q(\tag[1][11] ), 
        .QN(n1158) );
  DFFRX1 \tag_reg[1][10]  ( .D(n3134), .CK(clk), .RN(n3766), .Q(\tag[1][10] ), 
        .QN(n1157) );
  DFFRX1 \tag_reg[1][9]  ( .D(n3135), .CK(clk), .RN(n3766), .Q(\tag[1][9] ), 
        .QN(n1156) );
  DFFRX1 \tag_reg[1][8]  ( .D(n3136), .CK(clk), .RN(n3766), .Q(\tag[1][8] ), 
        .QN(n1155) );
  DFFRX1 \tag_reg[1][7]  ( .D(n3137), .CK(clk), .RN(n3766), .QN(n1154) );
  DFFRX1 \tag_reg[1][6]  ( .D(n3138), .CK(clk), .RN(n3766), .QN(n1153) );
  DFFRX1 \tag_reg[1][5]  ( .D(n3139), .CK(clk), .RN(n3766), .QN(n1152) );
  DFFRX1 \tag_reg[1][4]  ( .D(n3140), .CK(clk), .RN(n3766), .QN(n1151) );
  DFFRX1 \tag_reg[1][3]  ( .D(n3141), .CK(clk), .RN(n3766), .Q(\tag[1][3] ), 
        .QN(n1150) );
  DFFRX1 \tag_reg[1][2]  ( .D(n3142), .CK(clk), .RN(n3766), .QN(n1149) );
  DFFRX1 \tag_reg[1][1]  ( .D(n3143), .CK(clk), .RN(n3765), .Q(\tag[1][1] ), 
        .QN(n1148) );
  DFFRX1 \tag_reg[1][0]  ( .D(n3144), .CK(clk), .RN(n3765), .Q(\tag[1][0] ), 
        .QN(n1147) );
  DFFRX1 \valid_reg[4]  ( .D(n1708), .CK(clk), .RN(n3774), .Q(valid[4]), .QN(
        n1699) );
  DFFRX1 \tag_reg[4][24]  ( .D(n3045), .CK(clk), .RN(n3774), .Q(\tag[4][24] ), 
        .QN(n1246) );
  DFFRX1 \tag_reg[4][23]  ( .D(n3046), .CK(clk), .RN(n3774), .Q(\tag[4][23] ), 
        .QN(n1245) );
  DFFRX1 \tag_reg[4][22]  ( .D(n3047), .CK(clk), .RN(n3774), .Q(\tag[4][22] ), 
        .QN(n1244) );
  DFFRX1 \tag_reg[4][21]  ( .D(n3048), .CK(clk), .RN(n3774), .Q(\tag[4][21] ), 
        .QN(n1243) );
  DFFRX1 \tag_reg[4][20]  ( .D(n3049), .CK(clk), .RN(n3774), .QN(n1242) );
  DFFRX1 \tag_reg[4][19]  ( .D(n3050), .CK(clk), .RN(n3773), .QN(n1241) );
  DFFRX1 \tag_reg[4][18]  ( .D(n3051), .CK(clk), .RN(n3773), .Q(\tag[4][18] ), 
        .QN(n1240) );
  DFFRX1 \tag_reg[4][17]  ( .D(n3052), .CK(clk), .RN(n3773), .QN(n1239) );
  DFFRX1 \tag_reg[4][16]  ( .D(n3053), .CK(clk), .RN(n3773), .Q(\tag[4][16] ), 
        .QN(n1238) );
  DFFRX1 \tag_reg[4][15]  ( .D(n3054), .CK(clk), .RN(n3773), .Q(\tag[4][15] ), 
        .QN(n1237) );
  DFFRX1 \tag_reg[4][14]  ( .D(n3055), .CK(clk), .RN(n3773), .Q(\tag[4][14] ), 
        .QN(n1236) );
  DFFRX1 \tag_reg[4][13]  ( .D(n3056), .CK(clk), .RN(n3773), .Q(\tag[4][13] ), 
        .QN(n1235) );
  DFFRX1 \tag_reg[4][12]  ( .D(n3057), .CK(clk), .RN(n3773), .Q(\tag[4][12] ), 
        .QN(n1234) );
  DFFRX1 \tag_reg[4][11]  ( .D(n3058), .CK(clk), .RN(n3773), .Q(\tag[4][11] ), 
        .QN(n1233) );
  DFFRX1 \tag_reg[4][10]  ( .D(n3059), .CK(clk), .RN(n3773), .Q(\tag[4][10] ), 
        .QN(n1232) );
  DFFRX1 \tag_reg[4][9]  ( .D(n3060), .CK(clk), .RN(n3773), .Q(\tag[4][9] ), 
        .QN(n1231) );
  DFFRX1 \tag_reg[4][8]  ( .D(n3061), .CK(clk), .RN(n3773), .Q(\tag[4][8] ), 
        .QN(n1230) );
  DFFRX1 \tag_reg[4][7]  ( .D(n3062), .CK(clk), .RN(n3772), .QN(n1229) );
  DFFRX1 \tag_reg[4][6]  ( .D(n3063), .CK(clk), .RN(n3772), .QN(n1228) );
  DFFRX1 \tag_reg[4][5]  ( .D(n3064), .CK(clk), .RN(n3772), .QN(n1227) );
  DFFRX1 \tag_reg[4][4]  ( .D(n3065), .CK(clk), .RN(n3772), .QN(n1226) );
  DFFRX1 \tag_reg[4][3]  ( .D(n3066), .CK(clk), .RN(n3772), .Q(\tag[4][3] ), 
        .QN(n1225) );
  DFFRX1 \tag_reg[4][2]  ( .D(n3067), .CK(clk), .RN(n3772), .QN(n1224) );
  DFFRX1 \tag_reg[4][1]  ( .D(n3068), .CK(clk), .RN(n3772), .Q(\tag[4][1] ), 
        .QN(n1223) );
  DFFRX1 \tag_reg[4][0]  ( .D(n3069), .CK(clk), .RN(n3772), .Q(\tag[4][0] ), 
        .QN(n1222) );
  DFFRX1 \valid_reg[0]  ( .D(n1704), .CK(clk), .RN(n3765), .Q(valid[0]), .QN(
        n1703) );
  DFFRX1 \tag_reg[0][24]  ( .D(n3145), .CK(clk), .RN(n3765), .Q(\tag[0][24] ), 
        .QN(n1146) );
  DFFRX1 \tag_reg[0][23]  ( .D(n3146), .CK(clk), .RN(n3765), .Q(\tag[0][23] ), 
        .QN(n1145) );
  DFFRX1 \tag_reg[0][22]  ( .D(n3147), .CK(clk), .RN(n3765), .Q(\tag[0][22] ), 
        .QN(n1144) );
  DFFRX1 \tag_reg[0][21]  ( .D(n3148), .CK(clk), .RN(n3765), .Q(\tag[0][21] ), 
        .QN(n1143) );
  DFFRX1 \tag_reg[0][20]  ( .D(n3149), .CK(clk), .RN(n3765), .QN(n1142) );
  DFFRX1 \tag_reg[0][19]  ( .D(n3150), .CK(clk), .RN(n3765), .QN(n1141) );
  DFFRX1 \tag_reg[0][18]  ( .D(n3151), .CK(clk), .RN(n3765), .Q(\tag[0][18] ), 
        .QN(n1140) );
  DFFRX1 \tag_reg[0][17]  ( .D(n3152), .CK(clk), .RN(n3765), .QN(n1139) );
  DFFRX1 \tag_reg[0][16]  ( .D(n3153), .CK(clk), .RN(n3765), .Q(\tag[0][16] ), 
        .QN(n1138) );
  DFFRX1 \tag_reg[0][15]  ( .D(n3154), .CK(clk), .RN(n3764), .Q(\tag[0][15] ), 
        .QN(n1137) );
  DFFRX1 \tag_reg[0][14]  ( .D(n3155), .CK(clk), .RN(n3764), .Q(\tag[0][14] ), 
        .QN(n1136) );
  DFFRX1 \tag_reg[0][13]  ( .D(n3156), .CK(clk), .RN(n3764), .Q(\tag[0][13] ), 
        .QN(n1135) );
  DFFRX1 \tag_reg[0][12]  ( .D(n3157), .CK(clk), .RN(n3764), .Q(\tag[0][12] ), 
        .QN(n1134) );
  DFFRX1 \tag_reg[0][11]  ( .D(n3158), .CK(clk), .RN(n3764), .Q(\tag[0][11] ), 
        .QN(n1133) );
  DFFRX1 \tag_reg[0][10]  ( .D(n3159), .CK(clk), .RN(n3764), .Q(\tag[0][10] ), 
        .QN(n1132) );
  DFFRX1 \tag_reg[0][9]  ( .D(n3160), .CK(clk), .RN(n3764), .Q(\tag[0][9] ), 
        .QN(n1131) );
  DFFRX1 \tag_reg[0][8]  ( .D(n3161), .CK(clk), .RN(n3764), .Q(\tag[0][8] ), 
        .QN(n1130) );
  DFFRX1 \tag_reg[0][7]  ( .D(n3162), .CK(clk), .RN(n3764), .QN(n1129) );
  DFFRX1 \tag_reg[0][6]  ( .D(n3163), .CK(clk), .RN(n3764), .QN(n1128) );
  DFFRX1 \tag_reg[0][5]  ( .D(n3164), .CK(clk), .RN(n3764), .QN(n1127) );
  DFFRX1 \tag_reg[0][4]  ( .D(n3165), .CK(clk), .RN(n3764), .QN(n1126) );
  DFFRX1 \tag_reg[0][3]  ( .D(n3166), .CK(clk), .RN(n3763), .Q(\tag[0][3] ), 
        .QN(n1125) );
  DFFRX1 \tag_reg[0][2]  ( .D(n3167), .CK(clk), .RN(n3763), .QN(n1124) );
  DFFRX1 \tag_reg[0][1]  ( .D(n3168), .CK(clk), .RN(n3763), .Q(\tag[0][1] ), 
        .QN(n1123) );
  DFFRX1 \tag_reg[0][0]  ( .D(n3169), .CK(clk), .RN(n3763), .Q(\tag[0][0] ), 
        .QN(n1122) );
  DFFRX1 \valid_reg[6]  ( .D(n1710), .CK(clk), .RN(n3778), .Q(valid[6]), .QN(
        n1697) );
  DFFRX1 \tag_reg[6][24]  ( .D(n2995), .CK(clk), .RN(n3778), .Q(\tag[6][24] ), 
        .QN(n1296) );
  DFFRX1 \tag_reg[6][23]  ( .D(n2996), .CK(clk), .RN(n3778), .Q(\tag[6][23] ), 
        .QN(n1295) );
  DFFRX1 \tag_reg[6][22]  ( .D(n2997), .CK(clk), .RN(n3778), .Q(\tag[6][22] ), 
        .QN(n1294) );
  DFFRX1 \tag_reg[6][21]  ( .D(n2998), .CK(clk), .RN(n3778), .Q(\tag[6][21] ), 
        .QN(n1293) );
  DFFRX1 \tag_reg[6][20]  ( .D(n2999), .CK(clk), .RN(n3778), .QN(n1292) );
  DFFRX1 \tag_reg[6][19]  ( .D(n3000), .CK(clk), .RN(n3778), .QN(n1291) );
  DFFRX1 \tag_reg[6][18]  ( .D(n3001), .CK(clk), .RN(n3778), .Q(\tag[6][18] ), 
        .QN(n1290) );
  DFFRX1 \tag_reg[6][17]  ( .D(n3002), .CK(clk), .RN(n3778), .QN(n1289) );
  DFFRX1 \tag_reg[6][16]  ( .D(n3003), .CK(clk), .RN(n3778), .Q(\tag[6][16] ), 
        .QN(n1288) );
  DFFRX1 \tag_reg[6][15]  ( .D(n3004), .CK(clk), .RN(n3777), .Q(\tag[6][15] ), 
        .QN(n1287) );
  DFFRX1 \tag_reg[6][14]  ( .D(n3005), .CK(clk), .RN(n3777), .Q(\tag[6][14] ), 
        .QN(n1286) );
  DFFRX1 \tag_reg[6][13]  ( .D(n3006), .CK(clk), .RN(n3777), .Q(\tag[6][13] ), 
        .QN(n1285) );
  DFFRX1 \tag_reg[6][12]  ( .D(n3007), .CK(clk), .RN(n3777), .Q(\tag[6][12] ), 
        .QN(n1284) );
  DFFRX1 \tag_reg[6][11]  ( .D(n3008), .CK(clk), .RN(n3777), .Q(\tag[6][11] ), 
        .QN(n1283) );
  DFFRX1 \tag_reg[6][10]  ( .D(n3009), .CK(clk), .RN(n3777), .Q(\tag[6][10] ), 
        .QN(n1282) );
  DFFRX1 \tag_reg[6][9]  ( .D(n3010), .CK(clk), .RN(n3777), .Q(\tag[6][9] ), 
        .QN(n1281) );
  DFFRX1 \tag_reg[6][8]  ( .D(n3011), .CK(clk), .RN(n3777), .Q(\tag[6][8] ), 
        .QN(n1280) );
  DFFRX1 \tag_reg[6][7]  ( .D(n3012), .CK(clk), .RN(n3777), .QN(n1279) );
  DFFRX1 \tag_reg[6][6]  ( .D(n3013), .CK(clk), .RN(n3777), .QN(n1278) );
  DFFRX1 \tag_reg[6][5]  ( .D(n3014), .CK(clk), .RN(n3777), .QN(n1277) );
  DFFRX1 \tag_reg[6][4]  ( .D(n3015), .CK(clk), .RN(n3777), .QN(n1276) );
  DFFRX1 \tag_reg[6][3]  ( .D(n3016), .CK(clk), .RN(n3776), .Q(\tag[6][3] ), 
        .QN(n1275) );
  DFFRX1 \tag_reg[6][2]  ( .D(n3017), .CK(clk), .RN(n3776), .QN(n1274) );
  DFFRX1 \tag_reg[6][1]  ( .D(n3018), .CK(clk), .RN(n3776), .Q(\tag[6][1] ), 
        .QN(n1273) );
  DFFRX1 \tag_reg[6][0]  ( .D(n3019), .CK(clk), .RN(n3776), .Q(\tag[6][0] ), 
        .QN(n1272) );
  DFFRX1 \valid_reg[2]  ( .D(n1706), .CK(clk), .RN(n3770), .Q(valid[2]), .QN(
        n1701) );
  DFFRX1 \tag_reg[2][24]  ( .D(n3095), .CK(clk), .RN(n3770), .Q(\tag[2][24] ), 
        .QN(n1196) );
  DFFRX1 \tag_reg[2][23]  ( .D(n3096), .CK(clk), .RN(n3769), .Q(\tag[2][23] ), 
        .QN(n1195) );
  DFFRX1 \tag_reg[2][22]  ( .D(n3097), .CK(clk), .RN(n3769), .Q(\tag[2][22] ), 
        .QN(n1194) );
  DFFRX1 \tag_reg[2][21]  ( .D(n3098), .CK(clk), .RN(n3769), .Q(\tag[2][21] ), 
        .QN(n1193) );
  DFFRX1 \tag_reg[2][20]  ( .D(n3099), .CK(clk), .RN(n3769), .QN(n1192) );
  DFFRX1 \tag_reg[2][19]  ( .D(n3100), .CK(clk), .RN(n3769), .QN(n1191) );
  DFFRX1 \tag_reg[2][18]  ( .D(n3101), .CK(clk), .RN(n3769), .Q(\tag[2][18] ), 
        .QN(n1190) );
  DFFRX1 \tag_reg[2][17]  ( .D(n3102), .CK(clk), .RN(n3769), .QN(n1189) );
  DFFRX1 \tag_reg[2][16]  ( .D(n3103), .CK(clk), .RN(n3769), .Q(\tag[2][16] ), 
        .QN(n1188) );
  DFFRX1 \tag_reg[2][15]  ( .D(n3104), .CK(clk), .RN(n3769), .Q(\tag[2][15] ), 
        .QN(n1187) );
  DFFRX1 \tag_reg[2][14]  ( .D(n3105), .CK(clk), .RN(n3769), .Q(\tag[2][14] ), 
        .QN(n1186) );
  DFFRX1 \tag_reg[2][13]  ( .D(n3106), .CK(clk), .RN(n3769), .Q(\tag[2][13] ), 
        .QN(n1185) );
  DFFRX1 \tag_reg[2][12]  ( .D(n3107), .CK(clk), .RN(n3769), .Q(\tag[2][12] ), 
        .QN(n1184) );
  DFFRX1 \tag_reg[2][11]  ( .D(n3108), .CK(clk), .RN(n3768), .Q(\tag[2][11] ), 
        .QN(n1183) );
  DFFRX1 \tag_reg[2][10]  ( .D(n3109), .CK(clk), .RN(n3768), .Q(\tag[2][10] ), 
        .QN(n1182) );
  DFFRX1 \tag_reg[2][9]  ( .D(n3110), .CK(clk), .RN(n3768), .Q(\tag[2][9] ), 
        .QN(n1181) );
  DFFRX1 \tag_reg[2][8]  ( .D(n3111), .CK(clk), .RN(n3768), .Q(\tag[2][8] ), 
        .QN(n1180) );
  DFFRX1 \tag_reg[2][7]  ( .D(n3112), .CK(clk), .RN(n3768), .QN(n1179) );
  DFFRX1 \tag_reg[2][6]  ( .D(n3113), .CK(clk), .RN(n3768), .QN(n1178) );
  DFFRX1 \tag_reg[2][5]  ( .D(n3114), .CK(clk), .RN(n3768), .QN(n1177) );
  DFFRX1 \tag_reg[2][4]  ( .D(n3115), .CK(clk), .RN(n3768), .QN(n1176) );
  DFFRX1 \tag_reg[2][3]  ( .D(n3116), .CK(clk), .RN(n3768), .Q(\tag[2][3] ), 
        .QN(n1175) );
  DFFRX1 \tag_reg[2][2]  ( .D(n3117), .CK(clk), .RN(n3768), .QN(n1174) );
  DFFRX1 \tag_reg[2][1]  ( .D(n3118), .CK(clk), .RN(n3768), .Q(\tag[2][1] ), 
        .QN(n1173) );
  DFFRX1 \tag_reg[2][0]  ( .D(n3119), .CK(clk), .RN(n3768), .Q(\tag[2][0] ), 
        .QN(n1172) );
  DFFRX1 from_state_2_reg ( .D(n3172), .CK(clk), .RN(n3237), .Q(n3235), .QN(
        n1713) );
  DFFRX1 \next_proc_wdata_reg[31]  ( .D(n2781), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[31]) );
  DFFRX1 \next_proc_wdata_reg[30]  ( .D(n2782), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[30]) );
  DFFRX1 \next_proc_wdata_reg[29]  ( .D(n2783), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[29]) );
  DFFRX1 \next_proc_wdata_reg[28]  ( .D(n2784), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[28]) );
  DFFRX1 \next_proc_wdata_reg[27]  ( .D(n2785), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[27]) );
  DFFRX1 \next_proc_wdata_reg[26]  ( .D(n2786), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[26]) );
  DFFRX1 \next_proc_wdata_reg[25]  ( .D(n2787), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[25]) );
  DFFRX1 \next_proc_wdata_reg[24]  ( .D(n2788), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[24]) );
  DFFRX1 \next_proc_wdata_reg[23]  ( .D(n2789), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[23]) );
  DFFRX1 \next_proc_wdata_reg[22]  ( .D(n2790), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[22]) );
  DFFRX1 \next_proc_wdata_reg[21]  ( .D(n2791), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[21]) );
  DFFRX1 \next_proc_wdata_reg[20]  ( .D(n2792), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[20]) );
  DFFRX1 \next_proc_wdata_reg[19]  ( .D(n2793), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[19]) );
  DFFRX1 \next_proc_wdata_reg[18]  ( .D(n2794), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[18]) );
  DFFRX1 \next_proc_wdata_reg[17]  ( .D(n2795), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[17]) );
  DFFRX1 \next_proc_wdata_reg[16]  ( .D(n2796), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[16]) );
  DFFRX1 \next_proc_wdata_reg[15]  ( .D(n2797), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[15]) );
  DFFRX1 \next_proc_wdata_reg[14]  ( .D(n2798), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[14]) );
  DFFRX1 \next_proc_wdata_reg[13]  ( .D(n2799), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[13]) );
  DFFRX1 \next_proc_wdata_reg[12]  ( .D(n2800), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[12]) );
  DFFRX1 \next_proc_wdata_reg[11]  ( .D(n2801), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[11]) );
  DFFRX1 \next_proc_wdata_reg[10]  ( .D(n2802), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[10]) );
  DFFRX1 \next_proc_wdata_reg[9]  ( .D(n2803), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[9]) );
  DFFRX1 \next_proc_wdata_reg[8]  ( .D(n2804), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[8]) );
  DFFRX1 \next_proc_wdata_reg[7]  ( .D(n2805), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[7]) );
  DFFRX1 \next_proc_wdata_reg[6]  ( .D(n2806), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[6]) );
  DFFRX1 \next_proc_wdata_reg[5]  ( .D(n2807), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[5]) );
  DFFRX1 \next_proc_wdata_reg[4]  ( .D(n2808), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[4]) );
  DFFRX1 \next_proc_wdata_reg[3]  ( .D(n2809), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[3]) );
  DFFRX1 \next_proc_wdata_reg[2]  ( .D(n2810), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[2]) );
  DFFRX1 \next_proc_wdata_reg[1]  ( .D(n2811), .CK(clk), .RN(n3237), .Q(
        next_proc_wdata[1]) );
  DFFRX1 \next_proc_wdata_reg[0]  ( .D(n2812), .CK(clk), .RN(n3238), .Q(
        next_proc_wdata[0]) );
  DFFRX1 rw_status_reg ( .D(n2780), .CK(clk), .RN(n3237), .Q(rw_status), .QN(
        n4307) );
  DFFRX1 \state_reg[1]  ( .D(n3171), .CK(clk), .RN(n3238), .Q(state[1]), .QN(
        n4306) );
  DFFRX1 \state_reg[0]  ( .D(n3170), .CK(clk), .RN(n3237), .Q(state[0]) );
  DFFRX1 \prev_mem_wdata_reg[7]  ( .D(n2961), .CK(clk), .RN(n3238), .Q(
        mem_wdata[7]) );
  DFFRX1 \prev_mem_wdata_reg[6]  ( .D(n2962), .CK(clk), .RN(n3237), .Q(
        mem_wdata[6]) );
  DFFRX1 \prev_mem_wdata_reg[5]  ( .D(n2963), .CK(clk), .RN(n3238), .Q(
        mem_wdata[5]) );
  DFFRX1 \prev_mem_wdata_reg[4]  ( .D(n2964), .CK(clk), .RN(n3237), .Q(
        mem_wdata[4]) );
  DFFRX1 \prev_mem_wdata_reg[3]  ( .D(n2965), .CK(clk), .RN(n3238), .Q(
        mem_wdata[3]) );
  DFFRX1 \prev_mem_wdata_reg[2]  ( .D(n2966), .CK(clk), .RN(n3237), .Q(
        mem_wdata[2]) );
  DFFRX1 \prev_mem_wdata_reg[1]  ( .D(n2967), .CK(clk), .RN(n3238), .Q(
        mem_wdata[1]) );
  DFFRX1 \prev_mem_wdata_reg[0]  ( .D(n2968), .CK(clk), .RN(n3237), .Q(
        mem_wdata[0]) );
  DFFRX1 \prev_mem_wdata_reg[31]  ( .D(n2937), .CK(clk), .RN(n3238), .Q(
        mem_wdata[31]) );
  DFFRX1 \prev_mem_wdata_reg[30]  ( .D(n2938), .CK(clk), .RN(n3237), .Q(
        mem_wdata[30]) );
  DFFRX1 \prev_mem_wdata_reg[29]  ( .D(n2939), .CK(clk), .RN(n3238), .Q(
        mem_wdata[29]) );
  DFFRX1 \prev_mem_wdata_reg[28]  ( .D(n2940), .CK(clk), .RN(n3237), .Q(
        mem_wdata[28]) );
  DFFRX1 \prev_mem_wdata_reg[27]  ( .D(n2941), .CK(clk), .RN(n3238), .Q(
        mem_wdata[27]) );
  DFFRX1 \prev_mem_wdata_reg[26]  ( .D(n2942), .CK(clk), .RN(n3237), .Q(
        mem_wdata[26]) );
  DFFRX1 \prev_mem_wdata_reg[25]  ( .D(n2943), .CK(clk), .RN(n3238), .Q(
        mem_wdata[25]) );
  DFFRX1 \prev_mem_wdata_reg[24]  ( .D(n2944), .CK(clk), .RN(n3237), .Q(
        mem_wdata[24]) );
  DFFRX1 \prev_mem_wdata_reg[23]  ( .D(n2945), .CK(clk), .RN(n3238), .Q(
        mem_wdata[23]) );
  DFFRX1 \prev_mem_wdata_reg[22]  ( .D(n2946), .CK(clk), .RN(n3237), .Q(
        mem_wdata[22]) );
  DFFRX1 \prev_mem_wdata_reg[21]  ( .D(n2947), .CK(clk), .RN(n3238), .Q(
        mem_wdata[21]) );
  DFFRX1 \prev_mem_wdata_reg[20]  ( .D(n2948), .CK(clk), .RN(n3237), .Q(
        mem_wdata[20]) );
  DFFRX1 \prev_mem_wdata_reg[19]  ( .D(n2949), .CK(clk), .RN(n3238), .Q(
        mem_wdata[19]) );
  DFFRX1 \prev_mem_wdata_reg[18]  ( .D(n2950), .CK(clk), .RN(n3237), .Q(
        mem_wdata[18]) );
  DFFRX1 \prev_mem_wdata_reg[17]  ( .D(n2951), .CK(clk), .RN(n3238), .Q(
        mem_wdata[17]) );
  DFFRX1 \prev_mem_wdata_reg[16]  ( .D(n2952), .CK(clk), .RN(n3237), .Q(
        mem_wdata[16]) );
  DFFRX1 \prev_mem_wdata_reg[15]  ( .D(n2953), .CK(clk), .RN(n3238), .Q(
        mem_wdata[15]) );
  DFFRX1 \prev_mem_wdata_reg[14]  ( .D(n2954), .CK(clk), .RN(n3237), .Q(
        mem_wdata[14]) );
  DFFRX1 \prev_mem_wdata_reg[13]  ( .D(n2955), .CK(clk), .RN(n3238), .Q(
        mem_wdata[13]) );
  DFFRX1 \prev_mem_wdata_reg[12]  ( .D(n2956), .CK(clk), .RN(n3237), .Q(
        mem_wdata[12]) );
  DFFRX1 \prev_mem_wdata_reg[11]  ( .D(n2957), .CK(clk), .RN(n3238), .Q(
        mem_wdata[11]) );
  DFFRX1 \prev_mem_wdata_reg[10]  ( .D(n2958), .CK(clk), .RN(n3237), .Q(
        mem_wdata[10]) );
  DFFRX1 \prev_mem_wdata_reg[9]  ( .D(n2959), .CK(clk), .RN(n3238), .Q(
        mem_wdata[9]) );
  DFFRX1 \prev_mem_wdata_reg[8]  ( .D(n2960), .CK(clk), .RN(n3237), .Q(
        mem_wdata[8]) );
  DFFRX1 \prev_mem_wdata_reg[127]  ( .D(n2841), .CK(clk), .RN(n3238), .Q(
        mem_wdata[127]) );
  DFFRX1 \prev_mem_wdata_reg[126]  ( .D(n2842), .CK(clk), .RN(n3237), .Q(
        mem_wdata[126]) );
  DFFRX1 \prev_mem_wdata_reg[125]  ( .D(n2843), .CK(clk), .RN(n3238), .Q(
        mem_wdata[125]) );
  DFFRX1 \prev_mem_wdata_reg[124]  ( .D(n2844), .CK(clk), .RN(n3237), .Q(
        mem_wdata[124]) );
  DFFRX1 \prev_mem_wdata_reg[123]  ( .D(n2845), .CK(clk), .RN(n3238), .Q(
        mem_wdata[123]) );
  DFFRX1 \prev_mem_wdata_reg[122]  ( .D(n2846), .CK(clk), .RN(n3237), .Q(
        mem_wdata[122]) );
  DFFRX1 \prev_mem_wdata_reg[121]  ( .D(n2847), .CK(clk), .RN(n3238), .Q(
        mem_wdata[121]) );
  DFFRX1 \prev_mem_wdata_reg[120]  ( .D(n2848), .CK(clk), .RN(n3237), .Q(
        mem_wdata[120]) );
  DFFRX1 \prev_mem_wdata_reg[119]  ( .D(n2849), .CK(clk), .RN(n3238), .Q(
        mem_wdata[119]) );
  DFFRX1 \prev_mem_wdata_reg[118]  ( .D(n2850), .CK(clk), .RN(n3237), .Q(
        mem_wdata[118]) );
  DFFRX1 \prev_mem_wdata_reg[117]  ( .D(n2851), .CK(clk), .RN(n3238), .Q(
        mem_wdata[117]) );
  DFFRX1 \prev_mem_wdata_reg[116]  ( .D(n2852), .CK(clk), .RN(n3237), .Q(
        mem_wdata[116]) );
  DFFRX1 \prev_mem_wdata_reg[115]  ( .D(n2853), .CK(clk), .RN(n3238), .Q(
        mem_wdata[115]) );
  DFFRX1 \prev_mem_wdata_reg[114]  ( .D(n2854), .CK(clk), .RN(n3237), .Q(
        mem_wdata[114]) );
  DFFRX1 \prev_mem_wdata_reg[113]  ( .D(n2855), .CK(clk), .RN(n3238), .Q(
        mem_wdata[113]) );
  DFFRX1 \prev_mem_wdata_reg[112]  ( .D(n2856), .CK(clk), .RN(n3237), .Q(
        mem_wdata[112]) );
  DFFRX1 \prev_mem_wdata_reg[111]  ( .D(n2857), .CK(clk), .RN(n3238), .Q(
        mem_wdata[111]) );
  DFFRX1 \prev_mem_wdata_reg[110]  ( .D(n2858), .CK(clk), .RN(n3237), .Q(
        mem_wdata[110]) );
  DFFRX1 \prev_mem_wdata_reg[109]  ( .D(n2859), .CK(clk), .RN(n3238), .Q(
        mem_wdata[109]) );
  DFFRX1 \prev_mem_wdata_reg[108]  ( .D(n2860), .CK(clk), .RN(n3237), .Q(
        mem_wdata[108]) );
  DFFRX1 \prev_mem_wdata_reg[107]  ( .D(n2861), .CK(clk), .RN(n3238), .Q(
        mem_wdata[107]) );
  DFFRX1 \prev_mem_wdata_reg[106]  ( .D(n2862), .CK(clk), .RN(n3237), .Q(
        mem_wdata[106]) );
  DFFRX1 \prev_mem_wdata_reg[105]  ( .D(n2863), .CK(clk), .RN(n3238), .Q(
        mem_wdata[105]) );
  DFFRX1 \prev_mem_wdata_reg[104]  ( .D(n2864), .CK(clk), .RN(n3237), .Q(
        mem_wdata[104]) );
  DFFRX1 \prev_mem_wdata_reg[103]  ( .D(n2865), .CK(clk), .RN(n3238), .Q(
        mem_wdata[103]) );
  DFFRX1 \prev_mem_wdata_reg[102]  ( .D(n2866), .CK(clk), .RN(n3237), .Q(
        mem_wdata[102]) );
  DFFRX1 \prev_mem_wdata_reg[101]  ( .D(n2867), .CK(clk), .RN(n3238), .Q(
        mem_wdata[101]) );
  DFFRX1 \prev_mem_wdata_reg[100]  ( .D(n2868), .CK(clk), .RN(n3237), .Q(
        mem_wdata[100]) );
  DFFRX1 \prev_mem_wdata_reg[99]  ( .D(n2869), .CK(clk), .RN(n3238), .Q(
        mem_wdata[99]) );
  DFFRX1 \prev_mem_wdata_reg[98]  ( .D(n2870), .CK(clk), .RN(n3237), .Q(
        mem_wdata[98]) );
  DFFRX1 \prev_mem_wdata_reg[97]  ( .D(n2871), .CK(clk), .RN(n3238), .Q(
        mem_wdata[97]) );
  DFFRX1 \prev_mem_wdata_reg[96]  ( .D(n2872), .CK(clk), .RN(n3237), .Q(
        mem_wdata[96]) );
  DFFRX1 \prev_mem_wdata_reg[95]  ( .D(n2873), .CK(clk), .RN(n3238), .Q(
        mem_wdata[95]) );
  DFFRX1 \prev_mem_wdata_reg[94]  ( .D(n2874), .CK(clk), .RN(n3237), .Q(
        mem_wdata[94]) );
  DFFRX1 \prev_mem_wdata_reg[93]  ( .D(n2875), .CK(clk), .RN(n3238), .Q(
        mem_wdata[93]) );
  DFFRX1 \prev_mem_wdata_reg[92]  ( .D(n2876), .CK(clk), .RN(n3237), .Q(
        mem_wdata[92]) );
  DFFRX1 \prev_mem_wdata_reg[91]  ( .D(n2877), .CK(clk), .RN(n3238), .Q(
        mem_wdata[91]) );
  DFFRX1 \prev_mem_wdata_reg[90]  ( .D(n2878), .CK(clk), .RN(n3237), .Q(
        mem_wdata[90]) );
  DFFRX1 \prev_mem_wdata_reg[89]  ( .D(n2879), .CK(clk), .RN(n3238), .Q(
        mem_wdata[89]) );
  DFFRX1 \prev_mem_wdata_reg[88]  ( .D(n2880), .CK(clk), .RN(n3237), .Q(
        mem_wdata[88]) );
  DFFRX1 \prev_mem_wdata_reg[87]  ( .D(n2881), .CK(clk), .RN(n3238), .Q(
        mem_wdata[87]) );
  DFFRX1 \prev_mem_wdata_reg[86]  ( .D(n2882), .CK(clk), .RN(n3237), .Q(
        mem_wdata[86]) );
  DFFRX1 \prev_mem_wdata_reg[85]  ( .D(n2883), .CK(clk), .RN(n3238), .Q(
        mem_wdata[85]) );
  DFFRX1 \prev_mem_wdata_reg[84]  ( .D(n2884), .CK(clk), .RN(n3237), .Q(
        mem_wdata[84]) );
  DFFRX1 \prev_mem_wdata_reg[83]  ( .D(n2885), .CK(clk), .RN(n3238), .Q(
        mem_wdata[83]) );
  DFFRX1 \prev_mem_wdata_reg[82]  ( .D(n2886), .CK(clk), .RN(n3237), .Q(
        mem_wdata[82]) );
  DFFRX1 \prev_mem_wdata_reg[81]  ( .D(n2887), .CK(clk), .RN(n3238), .Q(
        mem_wdata[81]) );
  DFFRX1 \prev_mem_wdata_reg[80]  ( .D(n2888), .CK(clk), .RN(n3237), .Q(
        mem_wdata[80]) );
  DFFRX1 \prev_mem_wdata_reg[79]  ( .D(n2889), .CK(clk), .RN(n3238), .Q(
        mem_wdata[79]) );
  DFFRX1 \prev_mem_wdata_reg[78]  ( .D(n2890), .CK(clk), .RN(n3237), .Q(
        mem_wdata[78]) );
  DFFRX1 \prev_mem_wdata_reg[77]  ( .D(n2891), .CK(clk), .RN(n3238), .Q(
        mem_wdata[77]) );
  DFFRX1 \prev_mem_wdata_reg[76]  ( .D(n2892), .CK(clk), .RN(n3237), .Q(
        mem_wdata[76]) );
  DFFRX1 \prev_mem_wdata_reg[75]  ( .D(n2893), .CK(clk), .RN(n3238), .Q(
        mem_wdata[75]) );
  DFFRX1 \prev_mem_wdata_reg[74]  ( .D(n2894), .CK(clk), .RN(n3237), .Q(
        mem_wdata[74]) );
  DFFRX1 \prev_mem_wdata_reg[73]  ( .D(n2895), .CK(clk), .RN(n3238), .Q(
        mem_wdata[73]) );
  DFFRX1 \prev_mem_wdata_reg[72]  ( .D(n2896), .CK(clk), .RN(n3237), .Q(
        mem_wdata[72]) );
  DFFRX1 \prev_mem_wdata_reg[71]  ( .D(n2897), .CK(clk), .RN(n3238), .Q(
        mem_wdata[71]) );
  DFFRX1 \prev_mem_wdata_reg[70]  ( .D(n2898), .CK(clk), .RN(n3237), .Q(
        mem_wdata[70]) );
  DFFRX1 \prev_mem_wdata_reg[69]  ( .D(n2899), .CK(clk), .RN(n3238), .Q(
        mem_wdata[69]) );
  DFFRX1 \prev_mem_wdata_reg[68]  ( .D(n2900), .CK(clk), .RN(n3237), .Q(
        mem_wdata[68]) );
  DFFRX1 \prev_mem_wdata_reg[67]  ( .D(n2901), .CK(clk), .RN(n3238), .Q(
        mem_wdata[67]) );
  DFFRX1 \prev_mem_wdata_reg[66]  ( .D(n2902), .CK(clk), .RN(n3237), .Q(
        mem_wdata[66]) );
  DFFRX1 \prev_mem_wdata_reg[65]  ( .D(n2903), .CK(clk), .RN(n3238), .Q(
        mem_wdata[65]) );
  DFFRX1 \prev_mem_wdata_reg[64]  ( .D(n2904), .CK(clk), .RN(n3237), .Q(
        mem_wdata[64]) );
  DFFRX1 \prev_mem_wdata_reg[63]  ( .D(n2905), .CK(clk), .RN(n3238), .Q(
        mem_wdata[63]) );
  DFFRX1 \prev_mem_wdata_reg[62]  ( .D(n2906), .CK(clk), .RN(n3237), .Q(
        mem_wdata[62]) );
  DFFRX1 \prev_mem_wdata_reg[61]  ( .D(n2907), .CK(clk), .RN(n3238), .Q(
        mem_wdata[61]) );
  DFFRX1 \prev_mem_wdata_reg[60]  ( .D(n2908), .CK(clk), .RN(n3237), .Q(
        mem_wdata[60]) );
  DFFRX1 \prev_mem_wdata_reg[59]  ( .D(n2909), .CK(clk), .RN(n3238), .Q(
        mem_wdata[59]) );
  DFFRX1 \prev_mem_wdata_reg[58]  ( .D(n2910), .CK(clk), .RN(n3237), .Q(
        mem_wdata[58]) );
  DFFRX1 \prev_mem_wdata_reg[57]  ( .D(n2911), .CK(clk), .RN(n3238), .Q(
        mem_wdata[57]) );
  DFFRX1 \prev_mem_wdata_reg[56]  ( .D(n2912), .CK(clk), .RN(n3237), .Q(
        mem_wdata[56]) );
  DFFRX1 \prev_mem_wdata_reg[55]  ( .D(n2913), .CK(clk), .RN(n3238), .Q(
        mem_wdata[55]) );
  DFFRX1 \prev_mem_wdata_reg[54]  ( .D(n2914), .CK(clk), .RN(n3237), .Q(
        mem_wdata[54]) );
  DFFRX1 \prev_mem_wdata_reg[53]  ( .D(n2915), .CK(clk), .RN(n3238), .Q(
        mem_wdata[53]) );
  DFFRX1 \prev_mem_wdata_reg[52]  ( .D(n2916), .CK(clk), .RN(n3237), .Q(
        mem_wdata[52]) );
  DFFRX1 \prev_mem_wdata_reg[51]  ( .D(n2917), .CK(clk), .RN(n3238), .Q(
        mem_wdata[51]) );
  DFFRX1 \prev_mem_wdata_reg[50]  ( .D(n2918), .CK(clk), .RN(n3237), .Q(
        mem_wdata[50]) );
  DFFRX1 \prev_mem_wdata_reg[49]  ( .D(n2919), .CK(clk), .RN(n3238), .Q(
        mem_wdata[49]) );
  DFFRX1 \prev_mem_wdata_reg[48]  ( .D(n2920), .CK(clk), .RN(n3237), .Q(
        mem_wdata[48]) );
  DFFRX1 \prev_mem_wdata_reg[47]  ( .D(n2921), .CK(clk), .RN(n3238), .Q(
        mem_wdata[47]) );
  DFFRX1 \prev_mem_wdata_reg[46]  ( .D(n2922), .CK(clk), .RN(n3237), .Q(
        mem_wdata[46]) );
  DFFRX1 \prev_mem_wdata_reg[45]  ( .D(n2923), .CK(clk), .RN(n3238), .Q(
        mem_wdata[45]) );
  DFFRX1 \prev_mem_wdata_reg[44]  ( .D(n2924), .CK(clk), .RN(n3237), .Q(
        mem_wdata[44]) );
  DFFRX1 \prev_mem_wdata_reg[43]  ( .D(n2925), .CK(clk), .RN(n3238), .Q(
        mem_wdata[43]) );
  DFFRX1 \prev_mem_wdata_reg[42]  ( .D(n2926), .CK(clk), .RN(n3237), .Q(
        mem_wdata[42]) );
  DFFRX1 \prev_mem_wdata_reg[41]  ( .D(n2927), .CK(clk), .RN(n3238), .Q(
        mem_wdata[41]) );
  DFFRX1 \prev_mem_wdata_reg[40]  ( .D(n2928), .CK(clk), .RN(n3237), .Q(
        mem_wdata[40]) );
  DFFRX1 \prev_mem_wdata_reg[39]  ( .D(n2929), .CK(clk), .RN(n3238), .Q(
        mem_wdata[39]) );
  DFFRX1 \prev_mem_wdata_reg[38]  ( .D(n2930), .CK(clk), .RN(n3237), .Q(
        mem_wdata[38]) );
  DFFRX1 \prev_mem_wdata_reg[37]  ( .D(n2931), .CK(clk), .RN(n3238), .Q(
        mem_wdata[37]) );
  DFFRX1 \prev_mem_wdata_reg[36]  ( .D(n2932), .CK(clk), .RN(n3237), .Q(
        mem_wdata[36]) );
  DFFRX1 \prev_mem_wdata_reg[35]  ( .D(n2933), .CK(clk), .RN(n3238), .Q(
        mem_wdata[35]) );
  DFFRX1 \prev_mem_wdata_reg[34]  ( .D(n2934), .CK(clk), .RN(n3237), .Q(
        mem_wdata[34]) );
  DFFRX1 \prev_mem_wdata_reg[33]  ( .D(n2935), .CK(clk), .RN(n3238), .Q(
        mem_wdata[33]) );
  DFFRX1 \prev_mem_wdata_reg[32]  ( .D(n2936), .CK(clk), .RN(n3237), .Q(
        mem_wdata[32]) );
  OAI21X1 U1866 ( .A0(n3255), .A1(n309), .B0(n3937), .Y(n330) );
  CLKBUFX8 U1867 ( .A(n346), .Y(n3186) );
  CLKBUFX8 U1868 ( .A(n338), .Y(n3190) );
  CLKBUFX8 U1869 ( .A(n354), .Y(n3187) );
  CLKBUFX8 U1870 ( .A(n322), .Y(n3188) );
  OAI21X1 U1871 ( .A0(n3254), .A1(n305), .B0(n3950), .Y(n324) );
  CLKBUFX8 U1872 ( .A(n332), .Y(n3194) );
  CLKBUFX8 U1873 ( .A(n348), .Y(n3191) );
  CLKBUFX8 U1874 ( .A(n340), .Y(n3195) );
  CLKBUFX8 U1875 ( .A(n356), .Y(n3192) );
  OAI21X1 U1876 ( .A0(n102), .A1(n315), .B0(n3898), .Y(n360) );
  CLKBUFX8 U1877 ( .A(n336), .Y(n3199) );
  CLKBUFX8 U1878 ( .A(n328), .Y(n3200) );
  CLKBUFX8 U1879 ( .A(n344), .Y(n3196) );
  CLKBUFX8 U1880 ( .A(n352), .Y(n3197) );
  CLKBUFX8 U1881 ( .A(n364), .Y(n3201) );
  BUFX8 U1882 ( .A(n3270), .Y(n4025) );
  BUFX8 U1883 ( .A(n366), .Y(n3202) );
  BUFX8 U1884 ( .A(n3271), .Y(n4014) );
  OAI222X4 U1885 ( .A0(n406), .A1(n3268), .B0(n4109), .B1(n4038), .C0(n3885), 
        .C1(n4240), .Y(n2429) );
  OAI21X1 U1886 ( .A0(n3256), .A1(n101), .B0(n3884), .Y(n3268) );
  CLKBUFX6 U1887 ( .A(n3259), .Y(n3173) );
  INVX3 U1888 ( .A(n358), .Y(n3174) );
  CLKINVX12 U1889 ( .A(n3174), .Y(n3175) );
  INVX3 U1890 ( .A(n326), .Y(n3176) );
  CLKINVX12 U1891 ( .A(n3176), .Y(n3177) );
  INVX3 U1892 ( .A(n334), .Y(n3178) );
  CLKINVX12 U1893 ( .A(n3178), .Y(n3179) );
  INVX3 U1894 ( .A(n342), .Y(n3180) );
  CLKINVX12 U1895 ( .A(n3180), .Y(n3181) );
  INVX3 U1896 ( .A(n350), .Y(n3182) );
  CLKINVX12 U1897 ( .A(n3182), .Y(n3183) );
  XNOR2X1 U1898 ( .A(N217), .B(proc_addr[19]), .Y(n390) );
  XNOR2X1 U1899 ( .A(N222), .B(proc_addr[14]), .Y(n392) );
  NAND3X1 U1900 ( .A(n398), .B(n399), .C(n400), .Y(n394) );
  XNOR2X1 U1901 ( .A(N220), .B(proc_addr[16]), .Y(n398) );
  XNOR2X1 U1902 ( .A(N221), .B(proc_addr[15]), .Y(n399) );
  XNOR2X1 U1903 ( .A(N218), .B(proc_addr[18]), .Y(n400) );
  XNOR2X1 U1904 ( .A(N230), .B(proc_addr[6]), .Y(n377) );
  CLKBUFX3 U1905 ( .A(n3597), .Y(n3599) );
  BUFX4 U1906 ( .A(n184), .Y(n3256) );
  BUFX12 U1907 ( .A(n4118), .Y(n3623) );
  CLKBUFX3 U1908 ( .A(n3627), .Y(n3634) );
  CLKBUFX3 U1909 ( .A(n4114), .Y(n3659) );
  CLKBUFX6 U1910 ( .A(n3600), .Y(n3605) );
  CLKBUFX3 U1911 ( .A(n3600), .Y(n3604) );
  NAND2X2 U1912 ( .A(n3911), .B(n3183), .Y(n351) );
  CLKBUFX6 U1913 ( .A(n3269), .Y(n4015) );
  CLKBUFX6 U1914 ( .A(n3273), .Y(n4016) );
  NAND2X2 U1915 ( .A(n3924), .B(n3181), .Y(n343) );
  CLKBUFX6 U1916 ( .A(n3272), .Y(n4026) );
  CLKBUFX6 U1917 ( .A(n3274), .Y(n4027) );
  NAND2X2 U1918 ( .A(n3937), .B(n3179), .Y(n335) );
  NAND2X2 U1919 ( .A(n3898), .B(n3175), .Y(n359) );
  NAND2X2 U1920 ( .A(n3950), .B(n3177), .Y(n327) );
  CLKINVX16 U1921 ( .A(N42), .Y(n4119) );
  CLKINVX1 U1922 ( .A(N43), .Y(n4117) );
  MXI2X1 U1923 ( .A(n3304), .B(n3305), .S0(n3657), .Y(N214) );
  CLKBUFX6 U1924 ( .A(n3266), .Y(n3184) );
  NAND2X6 U1925 ( .A(n3860), .B(n4016), .Y(n3265) );
  NAND2X6 U1926 ( .A(n3860), .B(n4015), .Y(n3261) );
  CLKBUFX6 U1927 ( .A(n3264), .Y(n3185) );
  CLKBUFX6 U1928 ( .A(n330), .Y(n3189) );
  CLKBUFX6 U1929 ( .A(n324), .Y(n3193) );
  CLKBUFX6 U1930 ( .A(n360), .Y(n3198) );
  INVX3 U1931 ( .A(N44), .Y(n4115) );
  CLKINVX1 U1932 ( .A(n4115), .Y(n4114) );
  CLKBUFX2 U1933 ( .A(n3623), .Y(n3598) );
  OAI22X1 U1934 ( .A0(proc_wdata[2]), .A1(n3809), .B0(next_proc_wdata[2]), 
        .B1(n3807), .Y(n3203) );
  OAI22X1 U1935 ( .A0(proc_wdata[3]), .A1(n3235), .B0(next_proc_wdata[3]), 
        .B1(n3807), .Y(n3204) );
  OAI22X1 U1936 ( .A0(proc_wdata[28]), .A1(n3810), .B0(next_proc_wdata[28]), 
        .B1(n3807), .Y(n3205) );
  OAI22X1 U1937 ( .A0(proc_wdata[29]), .A1(n3811), .B0(next_proc_wdata[29]), 
        .B1(n3807), .Y(n3206) );
  OAI22X1 U1938 ( .A0(proc_wdata[30]), .A1(n3235), .B0(next_proc_wdata[30]), 
        .B1(n3807), .Y(n3207) );
  OAI22X1 U1939 ( .A0(proc_wdata[31]), .A1(n3810), .B0(next_proc_wdata[31]), 
        .B1(n3807), .Y(n3208) );
  BUFX8 U1940 ( .A(n3267), .Y(n4042) );
  OAI22X2 U1941 ( .A0(proc_wdata[24]), .A1(n3810), .B0(next_proc_wdata[24]), 
        .B1(n3808), .Y(n3209) );
  OAI22X1 U1942 ( .A0(proc_wdata[4]), .A1(n3810), .B0(next_proc_wdata[4]), 
        .B1(n3807), .Y(n3210) );
  OAI22X1 U1943 ( .A0(proc_wdata[5]), .A1(n3810), .B0(next_proc_wdata[5]), 
        .B1(n3807), .Y(n3211) );
  OAI22X1 U1944 ( .A0(proc_wdata[6]), .A1(n3810), .B0(next_proc_wdata[6]), 
        .B1(n3808), .Y(n3212) );
  OAI22X1 U1945 ( .A0(proc_wdata[7]), .A1(n3810), .B0(next_proc_wdata[7]), 
        .B1(n3808), .Y(n3213) );
  OAI22X1 U1946 ( .A0(proc_wdata[25]), .A1(n3809), .B0(next_proc_wdata[25]), 
        .B1(n3807), .Y(n3214) );
  OAI22X1 U1947 ( .A0(proc_wdata[26]), .A1(n3809), .B0(next_proc_wdata[26]), 
        .B1(n3807), .Y(n3215) );
  OAI22X1 U1948 ( .A0(proc_wdata[27]), .A1(n3809), .B0(next_proc_wdata[27]), 
        .B1(n3807), .Y(n3216) );
  OAI22X1 U1949 ( .A0(proc_wdata[0]), .A1(n3810), .B0(next_proc_wdata[0]), 
        .B1(n3808), .Y(n3217) );
  OAI22X1 U1950 ( .A0(proc_wdata[1]), .A1(n3810), .B0(next_proc_wdata[1]), 
        .B1(n3807), .Y(n3218) );
  OAI22X1 U1951 ( .A0(proc_wdata[8]), .A1(n3809), .B0(next_proc_wdata[8]), 
        .B1(n3808), .Y(n3219) );
  OAI22X1 U1952 ( .A0(proc_wdata[9]), .A1(n3809), .B0(next_proc_wdata[9]), 
        .B1(n3808), .Y(n3220) );
  OAI22X1 U1953 ( .A0(proc_wdata[10]), .A1(n3810), .B0(next_proc_wdata[10]), 
        .B1(n3808), .Y(n3221) );
  OAI22X1 U1954 ( .A0(proc_wdata[11]), .A1(n3810), .B0(next_proc_wdata[11]), 
        .B1(n3808), .Y(n3222) );
  OAI22X1 U1955 ( .A0(proc_wdata[12]), .A1(n3810), .B0(next_proc_wdata[12]), 
        .B1(n3808), .Y(n3223) );
  OAI22X1 U1956 ( .A0(proc_wdata[13]), .A1(n3235), .B0(next_proc_wdata[13]), 
        .B1(n3808), .Y(n3224) );
  OAI22X1 U1957 ( .A0(proc_wdata[14]), .A1(n3810), .B0(next_proc_wdata[14]), 
        .B1(n3808), .Y(n3225) );
  OAI22X1 U1958 ( .A0(proc_wdata[15]), .A1(n3811), .B0(next_proc_wdata[15]), 
        .B1(n3808), .Y(n3226) );
  OAI22X1 U1959 ( .A0(proc_wdata[16]), .A1(n3810), .B0(next_proc_wdata[16]), 
        .B1(n3808), .Y(n3227) );
  OAI22X1 U1960 ( .A0(proc_wdata[17]), .A1(n3811), .B0(next_proc_wdata[17]), 
        .B1(n3808), .Y(n3228) );
  OAI22X1 U1961 ( .A0(proc_wdata[18]), .A1(n3811), .B0(next_proc_wdata[18]), 
        .B1(n3808), .Y(n3229) );
  OAI22X1 U1962 ( .A0(proc_wdata[19]), .A1(n3235), .B0(next_proc_wdata[19]), 
        .B1(n3808), .Y(n3230) );
  OAI22X1 U1963 ( .A0(proc_wdata[20]), .A1(n3810), .B0(next_proc_wdata[20]), 
        .B1(n3808), .Y(n3231) );
  OAI22X1 U1964 ( .A0(proc_wdata[21]), .A1(n3810), .B0(next_proc_wdata[21]), 
        .B1(n3807), .Y(n3232) );
  OAI22X1 U1965 ( .A0(proc_wdata[22]), .A1(n3810), .B0(next_proc_wdata[22]), 
        .B1(n1713), .Y(n3233) );
  OAI22X1 U1966 ( .A0(proc_wdata[23]), .A1(n3235), .B0(next_proc_wdata[23]), 
        .B1(n3808), .Y(n3234) );
  NAND3XL U1967 ( .A(n265), .B(n199), .C(N233), .Y(n267) );
  CLKBUFX2 U1968 ( .A(n3656), .Y(n3626) );
  NAND2X2 U1969 ( .A(n3884), .B(n3202), .Y(n367) );
  NAND2X2 U1970 ( .A(n3898), .B(n3192), .Y(n357) );
  NAND2X2 U1971 ( .A(n3911), .B(n3191), .Y(n349) );
  NAND2X2 U1972 ( .A(n3924), .B(n3195), .Y(n341) );
  NAND2X2 U1973 ( .A(n3937), .B(n3194), .Y(n333) );
  NAND2X2 U1974 ( .A(n3950), .B(n3193), .Y(n325) );
  NAND2X2 U1975 ( .A(n3884), .B(n3201), .Y(n365) );
  NAND2X2 U1976 ( .A(n3898), .B(n3187), .Y(n355) );
  NAND2X2 U1977 ( .A(n3911), .B(n3186), .Y(n347) );
  NAND2X2 U1978 ( .A(n3924), .B(n3190), .Y(n339) );
  NAND2X2 U1979 ( .A(n3937), .B(n3189), .Y(n331) );
  NAND2X2 U1980 ( .A(n3950), .B(n3188), .Y(n323) );
  NAND2X2 U1981 ( .A(n3898), .B(n3198), .Y(n361) );
  NAND2X2 U1982 ( .A(n3911), .B(n3197), .Y(n353) );
  NAND2X2 U1983 ( .A(n3924), .B(n3196), .Y(n345) );
  NAND2X2 U1984 ( .A(n3937), .B(n3199), .Y(n337) );
  NAND2X2 U1985 ( .A(n3950), .B(n3200), .Y(n329) );
  NAND2X1 U1986 ( .A(n3860), .B(n4014), .Y(n3262) );
  NAND2X1 U1987 ( .A(n3872), .B(n4025), .Y(n3263) );
  NAND2X1 U1988 ( .A(n3872), .B(n4026), .Y(n3264) );
  NAND2X1 U1989 ( .A(n3872), .B(n4027), .Y(n3266) );
  NAND2X1 U1990 ( .A(n3860), .B(n4009), .Y(n3257) );
  NAND2X1 U1991 ( .A(n3872), .B(n4020), .Y(n3258) );
  NAND2X1 U1992 ( .A(n3884), .B(n4042), .Y(n3259) );
  OAI21XL U1993 ( .A0(n3256), .A1(n315), .B0(n3898), .Y(n358) );
  OAI21XL U1994 ( .A0(n3256), .A1(n313), .B0(n3911), .Y(n350) );
  OAI21XL U1995 ( .A0(n3256), .A1(n311), .B0(n3924), .Y(n342) );
  OAI21XL U1996 ( .A0(n3256), .A1(n309), .B0(n3937), .Y(n334) );
  OAI21XL U1997 ( .A0(n3256), .A1(n305), .B0(n3950), .Y(n326) );
  OAI21XL U1998 ( .A0(n3254), .A1(n315), .B0(n3898), .Y(n356) );
  OAI21XL U1999 ( .A0(n3254), .A1(n313), .B0(n3911), .Y(n348) );
  OAI21XL U2000 ( .A0(n3254), .A1(n311), .B0(n3924), .Y(n340) );
  OAI21XL U2001 ( .A0(n3254), .A1(n309), .B0(n3937), .Y(n332) );
  OAI21XL U2002 ( .A0(n3255), .A1(n315), .B0(n3898), .Y(n354) );
  OAI21XL U2003 ( .A0(n3255), .A1(n313), .B0(n3911), .Y(n346) );
  OAI21XL U2004 ( .A0(n3255), .A1(n311), .B0(n3924), .Y(n338) );
  OAI21XL U2005 ( .A0(n3255), .A1(n305), .B0(n3950), .Y(n322) );
  OAI21XL U2006 ( .A0(n102), .A1(n313), .B0(n3911), .Y(n352) );
  OAI21XL U2007 ( .A0(n102), .A1(n311), .B0(n3924), .Y(n344) );
  OAI21XL U2008 ( .A0(n102), .A1(n309), .B0(n3937), .Y(n336) );
  OAI21XL U2009 ( .A0(n102), .A1(n305), .B0(n3950), .Y(n328) );
  OAI21XL U2010 ( .A0(n101), .A1(n3254), .B0(n3884), .Y(n366) );
  OAI21XL U2011 ( .A0(n101), .A1(n3255), .B0(n3884), .Y(n364) );
  CLKINVX1 U2012 ( .A(n3251), .Y(N230) );
  NAND2X2 U2013 ( .A(n3249), .B(n3250), .Y(n3251) );
  INVX3 U2014 ( .A(n4120), .Y(n3236) );
  INVX16 U2015 ( .A(n3236), .Y(n3237) );
  INVX16 U2016 ( .A(n3236), .Y(n3238) );
  OR2XL U2017 ( .A(n403), .B(n4112), .Y(n3239) );
  OR2XL U2018 ( .A(n4109), .B(n4032), .Y(n3240) );
  OR2X1 U2019 ( .A(n3885), .B(n4243), .Y(n3241) );
  NAND3X1 U2020 ( .A(n3239), .B(n3240), .C(n3241), .Y(n2432) );
  OR2XL U2021 ( .A(n401), .B(n4112), .Y(n3242) );
  OR2XL U2022 ( .A(n4109), .B(n4028), .Y(n3243) );
  OR2X1 U2023 ( .A(n3884), .B(n4245), .Y(n3244) );
  NAND3X1 U2024 ( .A(n3242), .B(n3243), .C(n3244), .Y(n2434) );
  NAND2X2 U2025 ( .A(n3308), .B(n3245), .Y(n3246) );
  NAND2X1 U2026 ( .A(n3309), .B(n3658), .Y(n3247) );
  NAND2X2 U2027 ( .A(n3246), .B(n3247), .Y(n3248) );
  INVXL U2028 ( .A(n3658), .Y(n3245) );
  INVX3 U2029 ( .A(n3248), .Y(N216) );
  MXI4XL U2030 ( .A(\tag[0][15] ), .B(\tag[1][15] ), .C(\tag[2][15] ), .D(
        \tag[3][15] ), .S0(n3603), .S1(n3632), .Y(n3308) );
  BUFX4 U2031 ( .A(N44), .Y(n3658) );
  INVX20 U2032 ( .A(n4119), .Y(n4118) );
  NAND2X2 U2033 ( .A(n3336), .B(n4115), .Y(n3249) );
  NAND2X2 U2034 ( .A(n3337), .B(n3659), .Y(n3250) );
  MXI4XL U2035 ( .A(\tag[0][1] ), .B(\tag[1][1] ), .C(\tag[2][1] ), .D(
        \tag[3][1] ), .S0(n3606), .S1(n3634), .Y(n3336) );
  MXI4XL U2036 ( .A(\tag[4][1] ), .B(\tag[5][1] ), .C(\tag[6][1] ), .D(
        \tag[7][1] ), .S0(n3606), .S1(n3634), .Y(n3337) );
  CLKBUFX6 U2037 ( .A(n3260), .Y(n4109) );
  NAND2X1 U2038 ( .A(n3884), .B(n4112), .Y(n3260) );
  XNOR2X1 U2039 ( .A(n4131), .B(N214), .Y(n382) );
  MXI2X2 U2040 ( .A(n3292), .B(n3293), .S0(n3657), .Y(N207) );
  CLKMX2X4 U2041 ( .A(n3252), .B(n3253), .S0(n3245), .Y(N211) );
  MXI4XL U2042 ( .A(n1242), .B(n1267), .C(n1292), .D(n1317), .S0(n3603), .S1(
        n3631), .Y(n3252) );
  MXI4XL U2043 ( .A(n1142), .B(n1167), .C(n1192), .D(n1217), .S0(n3603), .S1(
        n3631), .Y(n3253) );
  NAND3X2 U2044 ( .A(n320), .B(n4174), .C(N46), .Y(n174) );
  BUFX12 U2045 ( .A(n174), .Y(n3254) );
  NAND3X2 U2046 ( .A(N45), .B(n320), .C(N46), .Y(n138) );
  BUFX12 U2047 ( .A(n138), .Y(n3255) );
  CLKBUFX3 U2048 ( .A(n3625), .Y(n3628) );
  CLKBUFX3 U2049 ( .A(n3629), .Y(n3630) );
  NAND3X1 U2050 ( .A(n320), .B(n4173), .C(N45), .Y(n184) );
  CLKBUFX2 U2051 ( .A(n3596), .Y(n3601) );
  CLKBUFX3 U2052 ( .A(n3629), .Y(n3631) );
  BUFX2 U2053 ( .A(N43), .Y(n3656) );
  NAND3X4 U2054 ( .A(n4174), .B(n4173), .C(n320), .Y(n102) );
  NOR2X1 U2055 ( .A(n198), .B(n4307), .Y(n3277) );
  MX4X1 U2056 ( .A(n1241), .B(n1266), .C(n1291), .D(n1316), .S0(n3603), .S1(
        n3631), .Y(n3301) );
  MX4X1 U2057 ( .A(n1141), .B(n1166), .C(n1191), .D(n1216), .S0(n3603), .S1(
        n3631), .Y(n3300) );
  CLKBUFX2 U2058 ( .A(n3627), .Y(n3635) );
  OAI21XL U2059 ( .A0(n101), .A1(n102), .B0(n3884), .Y(n3267) );
  INVXL U2060 ( .A(n261), .Y(n4122) );
  INVX3 U2061 ( .A(n3281), .Y(n4000) );
  NOR4X2 U2062 ( .A(n372), .B(n373), .C(n374), .D(n375), .Y(n371) );
  OAI21XL U2063 ( .A0(n3254), .A1(n190), .B0(n3860), .Y(n3269) );
  OAI21XL U2064 ( .A0(n3256), .A1(n139), .B0(n3872), .Y(n3270) );
  OAI21XL U2065 ( .A0(n3256), .A1(n190), .B0(n3860), .Y(n3271) );
  CLKINVX1 U2066 ( .A(n4117), .Y(n4116) );
  OAI21XL U2067 ( .A0(n139), .A1(n3254), .B0(n3872), .Y(n3272) );
  OAI21XL U2068 ( .A0(n3255), .A1(n190), .B0(n3860), .Y(n3273) );
  OAI21XL U2069 ( .A0(n3255), .A1(n139), .B0(n3872), .Y(n3274) );
  NAND3X1 U2070 ( .A(n4117), .B(n4115), .C(n4118), .Y(n139) );
  AOI21X1 U2071 ( .A0(n4172), .A1(n258), .B0(n260), .Y(n205) );
  NAND3X1 U2072 ( .A(n4117), .B(n4115), .C(n4119), .Y(n190) );
  CLKINVX1 U2073 ( .A(n4174), .Y(n3285) );
  NAND2X1 U2074 ( .A(n303), .B(n3810), .Y(n198) );
  NAND4X2 U2075 ( .A(n390), .B(n391), .C(n392), .D(n393), .Y(n386) );
  XNOR2X4 U2076 ( .A(N216), .B(proc_addr[20]), .Y(n391) );
  XNOR2X2 U2077 ( .A(N212), .B(proc_addr[24]), .Y(n393) );
  MX4XL U2078 ( .A(n1127), .B(n1152), .C(n1177), .D(n1202), .S0(n3605), .S1(
        n3633), .Y(n3328) );
  MX4XL U2079 ( .A(n1227), .B(n1252), .C(n1277), .D(n1302), .S0(n3605), .S1(
        n3633), .Y(n3329) );
  MX4XL U2080 ( .A(n1128), .B(n1153), .C(n1178), .D(n1203), .S0(n3605), .S1(
        n3633), .Y(n3326) );
  MX4XL U2081 ( .A(n1228), .B(n1253), .C(n1278), .D(n1303), .S0(n3605), .S1(
        n3633), .Y(n3327) );
  MX4XL U2082 ( .A(n1124), .B(n1149), .C(n1174), .D(n1199), .S0(n3605), .S1(
        n3634), .Y(n3334) );
  MX4XL U2083 ( .A(n1224), .B(n1249), .C(n1274), .D(n1299), .S0(n3605), .S1(
        n3634), .Y(n3335) );
  MX4XL U2084 ( .A(n1126), .B(n1151), .C(n1176), .D(n1201), .S0(n3605), .S1(
        n3633), .Y(n3330) );
  MX4XL U2085 ( .A(n1226), .B(n1251), .C(n1276), .D(n1301), .S0(n3605), .S1(
        n3633), .Y(n3331) );
  MX4XL U2086 ( .A(n1139), .B(n1164), .C(n1189), .D(n1214), .S0(n3603), .S1(
        n3631), .Y(n3304) );
  MX4XL U2087 ( .A(n1239), .B(n1264), .C(n1289), .D(n1314), .S0(n3603), .S1(
        n3631), .Y(n3305) );
  MX4XL U2088 ( .A(n1129), .B(n1154), .C(n1179), .D(n1204), .S0(n3605), .S1(
        n3633), .Y(n3324) );
  MX4XL U2089 ( .A(n1229), .B(n1254), .C(n1279), .D(n1304), .S0(n3605), .S1(
        n3633), .Y(n3325) );
  INVXL U2090 ( .A(N229), .Y(n4150) );
  INVXL U2091 ( .A(N228), .Y(n4151) );
  INVXL U2092 ( .A(N227), .Y(n4152) );
  INVXL U2093 ( .A(N226), .Y(n4153) );
  INVXL U2094 ( .A(N225), .Y(n4154) );
  INVXL U2095 ( .A(N224), .Y(n4155) );
  INVXL U2096 ( .A(N223), .Y(n4156) );
  INVXL U2097 ( .A(N222), .Y(n4157) );
  INVXL U2098 ( .A(N221), .Y(n4158) );
  INVXL U2099 ( .A(N220), .Y(n4159) );
  INVXL U2100 ( .A(N219), .Y(n4160) );
  INVXL U2101 ( .A(N218), .Y(n4161) );
  INVXL U2102 ( .A(N217), .Y(n4162) );
  INVXL U2103 ( .A(N215), .Y(n4163) );
  INVXL U2104 ( .A(N214), .Y(n4164) );
  INVXL U2105 ( .A(N213), .Y(n4165) );
  INVXL U2106 ( .A(N212), .Y(n4166) );
  INVXL U2107 ( .A(N211), .Y(n4167) );
  INVXL U2108 ( .A(N210), .Y(n4168) );
  INVXL U2109 ( .A(N209), .Y(n4169) );
  INVXL U2110 ( .A(N208), .Y(n4170) );
  INVXL U2111 ( .A(N207), .Y(n4171) );
  INVXL U2112 ( .A(N231), .Y(n4149) );
  CLKBUFX3 U2113 ( .A(n272), .Y(n3667) );
  MXI4XL U2114 ( .A(valid[4]), .B(valid[5]), .C(valid[6]), .D(valid[7]), .S0(
        n3602), .S1(n3630), .Y(n3291) );
  MXI4XL U2115 ( .A(valid[0]), .B(valid[1]), .C(valid[2]), .D(valid[3]), .S0(
        n3602), .S1(n3630), .Y(n3290) );
  MX2X1 U2116 ( .A(n3283), .B(n3284), .S0(n3657), .Y(N233) );
  MX4XL U2117 ( .A(dirty[0]), .B(dirty[1]), .C(dirty[2]), .D(dirty[3]), .S0(
        n3602), .S1(n3630), .Y(n3283) );
  MX4XL U2118 ( .A(dirty[4]), .B(dirty[5]), .C(dirty[6]), .D(dirty[7]), .S0(
        n4118), .S1(n3630), .Y(n3284) );
  CLKINVX1 U2119 ( .A(N46), .Y(n4173) );
  MXI2XL U2120 ( .A(n3354), .B(n3355), .S0(n3659), .Y(N54) );
  MXI2XL U2121 ( .A(n3352), .B(n3353), .S0(n3659), .Y(N53) );
  MXI2XL U2122 ( .A(n3350), .B(n3351), .S0(n3659), .Y(N52) );
  MXI2XL U2123 ( .A(n3348), .B(n3349), .S0(n3659), .Y(N51) );
  MXI4XL U2124 ( .A(\block[4][3][27] ), .B(\block[5][3][27] ), .C(
        \block[6][3][27] ), .D(\block[7][3][27] ), .S0(n3606), .S1(n3635), .Y(
        n3349) );
  MXI2XL U2125 ( .A(n3346), .B(n3347), .S0(n3659), .Y(N50) );
  MXI4XL U2126 ( .A(\block[0][3][28] ), .B(\block[1][3][28] ), .C(
        \block[2][3][28] ), .D(\block[3][3][28] ), .S0(n3606), .S1(n3635), .Y(
        n3346) );
  MXI4XL U2127 ( .A(\block[4][3][28] ), .B(\block[5][3][28] ), .C(
        \block[6][3][28] ), .D(\block[7][3][28] ), .S0(n3606), .S1(n3635), .Y(
        n3347) );
  MXI2XL U2128 ( .A(n3344), .B(n3345), .S0(n3659), .Y(N49) );
  MXI4XL U2129 ( .A(\block[0][3][29] ), .B(\block[1][3][29] ), .C(
        \block[2][3][29] ), .D(\block[3][3][29] ), .S0(n4118), .S1(n3635), .Y(
        n3344) );
  MXI4XL U2130 ( .A(\block[4][3][29] ), .B(\block[5][3][29] ), .C(
        \block[6][3][29] ), .D(\block[7][3][29] ), .S0(n3606), .S1(n3635), .Y(
        n3345) );
  MXI2XL U2131 ( .A(n3342), .B(n3343), .S0(n3659), .Y(N48) );
  MXI4XL U2132 ( .A(\block[0][3][30] ), .B(\block[1][3][30] ), .C(
        \block[2][3][30] ), .D(\block[3][3][30] ), .S0(n3623), .S1(n3634), .Y(
        n3342) );
  MXI4XL U2133 ( .A(\block[4][3][30] ), .B(\block[5][3][30] ), .C(
        \block[6][3][30] ), .D(\block[7][3][30] ), .S0(n3606), .S1(n3634), .Y(
        n3343) );
  MXI2XL U2134 ( .A(n3340), .B(n3341), .S0(n3659), .Y(N47) );
  MXI4XL U2135 ( .A(\block[0][3][31] ), .B(\block[1][3][31] ), .C(
        \block[2][3][31] ), .D(\block[3][3][31] ), .S0(n3623), .S1(n3634), .Y(
        n3340) );
  MXI4XL U2136 ( .A(\block[4][3][31] ), .B(\block[5][3][31] ), .C(
        \block[6][3][31] ), .D(\block[7][3][31] ), .S0(n3606), .S1(n3634), .Y(
        n3341) );
  NOR2BX1 U2137 ( .AN(mem_ready), .B(n290), .Y(n260) );
  OAI31XL U2138 ( .A0(n3809), .A1(proc_write), .A2(proc_read), .B0(n303), .Y(
        n295) );
  NAND2X1 U2139 ( .A(state[0]), .B(n4306), .Y(n290) );
  CLKINVX1 U2140 ( .A(N45), .Y(n4174) );
  CLKINVX1 U2141 ( .A(proc_reset), .Y(n4120) );
  INVX1 U2142 ( .A(n4119), .Y(n3275) );
  NOR2X8 U2143 ( .A(n199), .B(n4000), .Y(n3276) );
  OR2X8 U2144 ( .A(n3276), .B(n3277), .Y(n320) );
  NAND4X4 U2145 ( .A(n368), .B(n369), .C(n370), .D(n371), .Y(n199) );
  AOI21XL U2146 ( .A0(n202), .A1(N233), .B0(n320), .Y(n308) );
  CLKBUFX3 U2147 ( .A(n3257), .Y(n4008) );
  CLKBUFX3 U2148 ( .A(n3257), .Y(n4007) );
  CLKBUFX3 U2149 ( .A(n3258), .Y(n4019) );
  CLKBUFX3 U2150 ( .A(n3258), .Y(n4018) );
  CLKBUFX3 U2151 ( .A(n3262), .Y(n4013) );
  CLKBUFX3 U2152 ( .A(n3262), .Y(n4012) );
  CLKBUFX3 U2153 ( .A(n3263), .Y(n4024) );
  CLKBUFX3 U2154 ( .A(n3263), .Y(n4023) );
  CLKBUFX3 U2155 ( .A(n3628), .Y(n3632) );
  CLKBUFX3 U2156 ( .A(n3628), .Y(n3633) );
  CLKBUFX3 U2157 ( .A(n3257), .Y(n4006) );
  CLKBUFX3 U2158 ( .A(n3258), .Y(n4017) );
  CLKBUFX3 U2159 ( .A(n3638), .Y(n3639) );
  CLKBUFX3 U2160 ( .A(n3626), .Y(n3654) );
  CLKBUFX3 U2161 ( .A(n3626), .Y(n3644) );
  CLKBUFX3 U2162 ( .A(n3636), .Y(n3648) );
  CLKBUFX3 U2163 ( .A(n3626), .Y(n3638) );
  CLKBUFX3 U2164 ( .A(n3626), .Y(n3653) );
  CLKBUFX3 U2165 ( .A(n3637), .Y(n3643) );
  CLKBUFX3 U2166 ( .A(n3649), .Y(n3647) );
  CLKBUFX3 U2167 ( .A(n3626), .Y(n3637) );
  CLKBUFX3 U2168 ( .A(n3626), .Y(n3652) );
  CLKBUFX3 U2169 ( .A(n3626), .Y(n3642) );
  CLKBUFX3 U2170 ( .A(n3626), .Y(n3646) );
  CLKBUFX3 U2171 ( .A(n3626), .Y(n3636) );
  CLKBUFX3 U2172 ( .A(n3626), .Y(n3651) );
  CLKBUFX3 U2173 ( .A(n3626), .Y(n3641) );
  CLKBUFX3 U2174 ( .A(n3635), .Y(n3650) );
  CLKBUFX3 U2175 ( .A(n3642), .Y(n3645) );
  CLKBUFX3 U2176 ( .A(n3626), .Y(n3649) );
  CLKBUFX3 U2177 ( .A(n3644), .Y(n3640) );
  CLKBUFX3 U2178 ( .A(n3599), .Y(n3606) );
  CLKBUFX3 U2179 ( .A(n3601), .Y(n3603) );
  CLKBUFX3 U2180 ( .A(n3601), .Y(n3602) );
  CLKBUFX3 U2181 ( .A(n361), .Y(n3817) );
  CLKBUFX3 U2182 ( .A(n361), .Y(n3816) );
  CLKBUFX3 U2183 ( .A(n353), .Y(n3825) );
  CLKBUFX3 U2184 ( .A(n353), .Y(n3824) );
  CLKBUFX3 U2185 ( .A(n345), .Y(n3833) );
  CLKBUFX3 U2186 ( .A(n345), .Y(n3832) );
  CLKBUFX3 U2187 ( .A(n337), .Y(n3841) );
  CLKBUFX3 U2188 ( .A(n337), .Y(n3840) );
  CLKBUFX3 U2189 ( .A(n329), .Y(n3849) );
  CLKBUFX3 U2190 ( .A(n329), .Y(n3848) );
  CLKBUFX3 U2191 ( .A(n3262), .Y(n4011) );
  CLKBUFX3 U2192 ( .A(n3263), .Y(n4022) );
  CLKBUFX3 U2193 ( .A(n3625), .Y(n3627) );
  INVX3 U2194 ( .A(n3867), .Y(n3860) );
  INVX3 U2195 ( .A(n3881), .Y(n3872) );
  INVX3 U2196 ( .A(n3906), .Y(n3898) );
  INVX3 U2197 ( .A(n3919), .Y(n3911) );
  INVX3 U2198 ( .A(n3932), .Y(n3924) );
  INVX3 U2199 ( .A(n3945), .Y(n3937) );
  INVX3 U2200 ( .A(n3958), .Y(n3950) );
  INVX3 U2201 ( .A(n3893), .Y(n3884) );
  INVX3 U2202 ( .A(n3969), .Y(n3965) );
  INVX3 U2203 ( .A(n3996), .Y(n3964) );
  INVX3 U2204 ( .A(n3971), .Y(n3963) );
  INVX3 U2205 ( .A(n3997), .Y(n3962) );
  INVX3 U2206 ( .A(n3997), .Y(n3961) );
  INVX3 U2207 ( .A(n3969), .Y(n3967) );
  INVX3 U2208 ( .A(n3970), .Y(n3966) );
  INVX3 U2209 ( .A(n3996), .Y(n3968) );
  CLKBUFX3 U2210 ( .A(n3664), .Y(n3660) );
  CLKBUFX3 U2211 ( .A(n3659), .Y(n3663) );
  CLKBUFX3 U2212 ( .A(n3663), .Y(n3662) );
  CLKBUFX3 U2213 ( .A(n3661), .Y(n3665) );
  CLKBUFX3 U2214 ( .A(n3659), .Y(n3664) );
  CLKBUFX3 U2215 ( .A(n3659), .Y(n3661) );
  CLKBUFX3 U2216 ( .A(n3598), .Y(n3618) );
  CLKBUFX3 U2217 ( .A(n3615), .Y(n3622) );
  CLKBUFX3 U2218 ( .A(n3598), .Y(n3610) );
  CLKBUFX3 U2219 ( .A(n3598), .Y(n3615) );
  CLKBUFX3 U2220 ( .A(n3607), .Y(n3621) );
  CLKBUFX3 U2221 ( .A(n3607), .Y(n3617) );
  CLKBUFX3 U2222 ( .A(n3598), .Y(n3614) );
  CLKBUFX3 U2223 ( .A(n3598), .Y(n3609) );
  CLKBUFX3 U2224 ( .A(n3607), .Y(n3620) );
  CLKBUFX3 U2225 ( .A(n3598), .Y(n3608) );
  CLKBUFX3 U2226 ( .A(n3598), .Y(n3613) );
  CLKBUFX3 U2227 ( .A(n3598), .Y(n3619) );
  CLKBUFX3 U2228 ( .A(n3598), .Y(n3616) );
  CLKBUFX3 U2229 ( .A(n3598), .Y(n3612) );
  CLKBUFX3 U2230 ( .A(n3599), .Y(n3607) );
  CLKBUFX3 U2231 ( .A(n3598), .Y(n3611) );
  INVX3 U2232 ( .A(n3905), .Y(n3900) );
  INVX3 U2233 ( .A(n3918), .Y(n3913) );
  INVX3 U2234 ( .A(n3931), .Y(n3926) );
  INVX3 U2235 ( .A(n3944), .Y(n3939) );
  INVX3 U2236 ( .A(n3957), .Y(n3952) );
  INVX3 U2237 ( .A(n3880), .Y(n3875) );
  INVX3 U2238 ( .A(n3905), .Y(n3901) );
  INVX3 U2239 ( .A(n3905), .Y(n3902) );
  INVX3 U2240 ( .A(n3918), .Y(n3914) );
  INVX3 U2241 ( .A(n3918), .Y(n3915) );
  INVX3 U2242 ( .A(n3931), .Y(n3927) );
  INVX3 U2243 ( .A(n3931), .Y(n3928) );
  INVX3 U2244 ( .A(n3944), .Y(n3940) );
  INVX3 U2245 ( .A(n3944), .Y(n3941) );
  INVX3 U2246 ( .A(n3957), .Y(n3953) );
  INVX3 U2247 ( .A(n3957), .Y(n3954) );
  INVX3 U2248 ( .A(n3866), .Y(n3862) );
  INVX3 U2249 ( .A(n3866), .Y(n3863) );
  INVX3 U2250 ( .A(n3907), .Y(n3903) );
  INVX3 U2251 ( .A(n3907), .Y(n3904) );
  INVX3 U2252 ( .A(n3920), .Y(n3916) );
  INVX3 U2253 ( .A(n3920), .Y(n3917) );
  INVX3 U2254 ( .A(n3933), .Y(n3929) );
  INVX3 U2255 ( .A(n3933), .Y(n3930) );
  INVX3 U2256 ( .A(n3946), .Y(n3942) );
  INVX3 U2257 ( .A(n3946), .Y(n3943) );
  INVX3 U2258 ( .A(n3959), .Y(n3955) );
  INVX3 U2259 ( .A(n3959), .Y(n3956) );
  INVX3 U2260 ( .A(n3868), .Y(n3864) );
  INVX3 U2261 ( .A(n3868), .Y(n3865) );
  INVX3 U2262 ( .A(n3907), .Y(n3899) );
  INVX3 U2263 ( .A(n3920), .Y(n3912) );
  INVX3 U2264 ( .A(n3933), .Y(n3925) );
  INVX3 U2265 ( .A(n3946), .Y(n3938) );
  INVX3 U2266 ( .A(n3959), .Y(n3951) );
  INVX3 U2267 ( .A(n3868), .Y(n3861) );
  INVX3 U2268 ( .A(n3870), .Y(n3873) );
  INVX3 U2269 ( .A(n3870), .Y(n3874) );
  INVX3 U2270 ( .A(n3880), .Y(n3876) );
  INVX3 U2271 ( .A(n3880), .Y(n3877) );
  INVX3 U2272 ( .A(n3892), .Y(n3885) );
  INVX3 U2273 ( .A(n3892), .Y(n3886) );
  INVX3 U2274 ( .A(n3892), .Y(n3887) );
  INVX3 U2275 ( .A(n3880), .Y(n3878) );
  INVX3 U2276 ( .A(n3880), .Y(n3879) );
  INVX3 U2277 ( .A(n3892), .Y(n3888) );
  INVX3 U2278 ( .A(n3892), .Y(n3889) );
  INVX3 U2279 ( .A(n3892), .Y(n3890) );
  INVX3 U2280 ( .A(n3868), .Y(n3858) );
  INVX3 U2281 ( .A(n3868), .Y(n3859) );
  INVX3 U2282 ( .A(n3880), .Y(n3871) );
  INVX3 U2283 ( .A(n3892), .Y(n3883) );
  INVX3 U2284 ( .A(n3907), .Y(n3897) );
  INVX3 U2285 ( .A(n3920), .Y(n3910) );
  INVX3 U2286 ( .A(n3933), .Y(n3923) );
  INVX3 U2287 ( .A(n3946), .Y(n3936) );
  INVX3 U2288 ( .A(n3959), .Y(n3949) );
  INVX3 U2289 ( .A(n3892), .Y(n3891) );
  CLKBUFX3 U2290 ( .A(N44), .Y(n3657) );
  CLKBUFX3 U2291 ( .A(n195), .Y(n4009) );
  CLKBUFX3 U2292 ( .A(n185), .Y(n4020) );
  CLKBUFX3 U2293 ( .A(n359), .Y(n3819) );
  CLKBUFX3 U2294 ( .A(n359), .Y(n3818) );
  CLKBUFX3 U2295 ( .A(n351), .Y(n3827) );
  CLKBUFX3 U2296 ( .A(n351), .Y(n3826) );
  CLKBUFX3 U2297 ( .A(n343), .Y(n3835) );
  CLKBUFX3 U2298 ( .A(n343), .Y(n3834) );
  CLKBUFX3 U2299 ( .A(n335), .Y(n3843) );
  CLKBUFX3 U2300 ( .A(n335), .Y(n3842) );
  CLKBUFX3 U2301 ( .A(n327), .Y(n3851) );
  CLKBUFX3 U2302 ( .A(n327), .Y(n3850) );
  CLKBUFX3 U2303 ( .A(n367), .Y(n3813) );
  CLKBUFX3 U2304 ( .A(n367), .Y(n3812) );
  CLKBUFX3 U2305 ( .A(n357), .Y(n3821) );
  CLKBUFX3 U2306 ( .A(n357), .Y(n3820) );
  CLKBUFX3 U2307 ( .A(n349), .Y(n3829) );
  CLKBUFX3 U2308 ( .A(n349), .Y(n3828) );
  CLKBUFX3 U2309 ( .A(n341), .Y(n3837) );
  CLKBUFX3 U2310 ( .A(n341), .Y(n3836) );
  CLKBUFX3 U2311 ( .A(n333), .Y(n3845) );
  CLKBUFX3 U2312 ( .A(n333), .Y(n3844) );
  CLKBUFX3 U2313 ( .A(n325), .Y(n3853) );
  CLKBUFX3 U2314 ( .A(n325), .Y(n3852) );
  CLKBUFX3 U2315 ( .A(n365), .Y(n3815) );
  CLKBUFX3 U2316 ( .A(n365), .Y(n3814) );
  CLKBUFX3 U2317 ( .A(n355), .Y(n3823) );
  CLKBUFX3 U2318 ( .A(n355), .Y(n3822) );
  CLKBUFX3 U2319 ( .A(n347), .Y(n3831) );
  CLKBUFX3 U2320 ( .A(n347), .Y(n3830) );
  CLKBUFX3 U2321 ( .A(n339), .Y(n3839) );
  CLKBUFX3 U2322 ( .A(n339), .Y(n3838) );
  CLKBUFX3 U2323 ( .A(n331), .Y(n3847) );
  CLKBUFX3 U2324 ( .A(n331), .Y(n3846) );
  CLKBUFX3 U2325 ( .A(n323), .Y(n3855) );
  CLKBUFX3 U2326 ( .A(n323), .Y(n3854) );
  CLKBUFX3 U2327 ( .A(n3656), .Y(n3625) );
  CLKBUFX3 U2328 ( .A(n3596), .Y(n3600) );
  CLKBUFX3 U2329 ( .A(n3856), .Y(n3867) );
  CLKBUFX3 U2330 ( .A(n3869), .Y(n3881) );
  CLKBUFX3 U2331 ( .A(n3882), .Y(n3893) );
  CLKBUFX3 U2332 ( .A(n3895), .Y(n3906) );
  CLKBUFX3 U2333 ( .A(n3908), .Y(n3919) );
  CLKBUFX3 U2334 ( .A(n3921), .Y(n3932) );
  CLKBUFX3 U2335 ( .A(n3934), .Y(n3945) );
  CLKBUFX3 U2336 ( .A(n3947), .Y(n3958) );
  CLKBUFX3 U2337 ( .A(n3960), .Y(n3971) );
  CLKBUFX3 U2338 ( .A(n3960), .Y(n3969) );
  CLKBUFX3 U2339 ( .A(n3960), .Y(n3970) );
  CLKBUFX3 U2340 ( .A(n4009), .Y(n4010) );
  CLKBUFX3 U2341 ( .A(n4020), .Y(n4021) );
  CLKBUFX3 U2342 ( .A(n3992), .Y(n3990) );
  CLKBUFX3 U2343 ( .A(n3992), .Y(n3989) );
  CLKBUFX3 U2344 ( .A(n3992), .Y(n3988) );
  CLKBUFX3 U2345 ( .A(n3993), .Y(n3987) );
  CLKBUFX3 U2346 ( .A(n3993), .Y(n3986) );
  CLKBUFX3 U2347 ( .A(n3993), .Y(n3985) );
  CLKBUFX3 U2348 ( .A(n3993), .Y(n3984) );
  CLKBUFX3 U2349 ( .A(n3994), .Y(n3983) );
  CLKBUFX3 U2350 ( .A(n3994), .Y(n3982) );
  CLKBUFX3 U2351 ( .A(n3994), .Y(n3981) );
  CLKBUFX3 U2352 ( .A(n3994), .Y(n3980) );
  CLKBUFX3 U2353 ( .A(n3995), .Y(n3979) );
  CLKBUFX3 U2354 ( .A(n3995), .Y(n3978) );
  CLKBUFX3 U2355 ( .A(n3995), .Y(n3977) );
  CLKBUFX3 U2356 ( .A(n3995), .Y(n3976) );
  CLKBUFX3 U2357 ( .A(n3996), .Y(n3975) );
  CLKBUFX3 U2358 ( .A(n3996), .Y(n3974) );
  CLKBUFX3 U2359 ( .A(n3996), .Y(n3973) );
  CLKBUFX3 U2360 ( .A(n3996), .Y(n3972) );
  CLKBUFX3 U2361 ( .A(n3992), .Y(n3991) );
  CLKBUFX3 U2362 ( .A(n3661), .Y(n3666) );
  CLKBUFX3 U2363 ( .A(n3856), .Y(n3868) );
  CLKBUFX3 U2364 ( .A(n3868), .Y(n3866) );
  CLKBUFX3 U2365 ( .A(n3881), .Y(n3880) );
  CLKBUFX3 U2366 ( .A(n3892), .Y(n3894) );
  CLKBUFX3 U2367 ( .A(n3882), .Y(n3892) );
  CLKBUFX3 U2368 ( .A(n3895), .Y(n3907) );
  CLKBUFX3 U2369 ( .A(n3907), .Y(n3905) );
  CLKBUFX3 U2370 ( .A(n3908), .Y(n3920) );
  CLKBUFX3 U2371 ( .A(n3920), .Y(n3918) );
  CLKBUFX3 U2372 ( .A(n3921), .Y(n3933) );
  CLKBUFX3 U2373 ( .A(n3933), .Y(n3931) );
  CLKBUFX3 U2374 ( .A(n3934), .Y(n3946) );
  CLKBUFX3 U2375 ( .A(n3946), .Y(n3944) );
  CLKBUFX3 U2376 ( .A(n3947), .Y(n3959) );
  CLKBUFX3 U2377 ( .A(n3959), .Y(n3957) );
  CLKBUFX3 U2378 ( .A(n3796), .Y(n3674) );
  CLKBUFX3 U2379 ( .A(n3796), .Y(n3675) );
  CLKBUFX3 U2380 ( .A(n3796), .Y(n3676) );
  CLKBUFX3 U2381 ( .A(n3796), .Y(n3677) );
  CLKBUFX3 U2382 ( .A(n3797), .Y(n3678) );
  CLKBUFX3 U2383 ( .A(n3797), .Y(n3679) );
  CLKBUFX3 U2384 ( .A(n3786), .Y(n3680) );
  CLKBUFX3 U2385 ( .A(n3785), .Y(n3681) );
  CLKBUFX3 U2386 ( .A(n3795), .Y(n3682) );
  CLKBUFX3 U2387 ( .A(n3795), .Y(n3683) );
  CLKBUFX3 U2388 ( .A(n3795), .Y(n3684) );
  CLKBUFX3 U2389 ( .A(n3795), .Y(n3685) );
  CLKBUFX3 U2390 ( .A(n3794), .Y(n3686) );
  CLKBUFX3 U2391 ( .A(n3794), .Y(n3687) );
  CLKBUFX3 U2392 ( .A(n3794), .Y(n3688) );
  CLKBUFX3 U2393 ( .A(n3794), .Y(n3689) );
  CLKBUFX3 U2394 ( .A(n3793), .Y(n3690) );
  CLKBUFX3 U2395 ( .A(n3793), .Y(n3691) );
  CLKBUFX3 U2396 ( .A(n3793), .Y(n3692) );
  CLKBUFX3 U2397 ( .A(n3793), .Y(n3693) );
  CLKBUFX3 U2398 ( .A(n3792), .Y(n3694) );
  CLKBUFX3 U2399 ( .A(n3792), .Y(n3695) );
  CLKBUFX3 U2400 ( .A(n3792), .Y(n3696) );
  CLKBUFX3 U2401 ( .A(n3792), .Y(n3697) );
  CLKBUFX3 U2402 ( .A(n3798), .Y(n3698) );
  CLKBUFX3 U2403 ( .A(n3798), .Y(n3699) );
  CLKBUFX3 U2404 ( .A(n3669), .Y(n3700) );
  CLKBUFX3 U2405 ( .A(n3787), .Y(n3701) );
  CLKBUFX3 U2406 ( .A(n3791), .Y(n3702) );
  CLKBUFX3 U2407 ( .A(n3791), .Y(n3703) );
  CLKBUFX3 U2408 ( .A(n3791), .Y(n3704) );
  CLKBUFX3 U2409 ( .A(n3791), .Y(n3705) );
  CLKBUFX3 U2410 ( .A(n3790), .Y(n3706) );
  CLKBUFX3 U2411 ( .A(n3790), .Y(n3707) );
  CLKBUFX3 U2412 ( .A(n3790), .Y(n3708) );
  CLKBUFX3 U2413 ( .A(n3790), .Y(n3709) );
  CLKBUFX3 U2414 ( .A(n3789), .Y(n3710) );
  CLKBUFX3 U2415 ( .A(n3789), .Y(n3711) );
  CLKBUFX3 U2416 ( .A(n3789), .Y(n3712) );
  CLKBUFX3 U2417 ( .A(n3789), .Y(n3713) );
  CLKBUFX3 U2418 ( .A(n3788), .Y(n3714) );
  CLKBUFX3 U2419 ( .A(n3788), .Y(n3715) );
  CLKBUFX3 U2420 ( .A(n3788), .Y(n3716) );
  CLKBUFX3 U2421 ( .A(n3788), .Y(n3717) );
  CLKBUFX3 U2422 ( .A(n3787), .Y(n3718) );
  CLKBUFX3 U2423 ( .A(n3787), .Y(n3719) );
  CLKBUFX3 U2424 ( .A(n3787), .Y(n3720) );
  CLKBUFX3 U2425 ( .A(n3787), .Y(n3721) );
  CLKBUFX3 U2426 ( .A(n3786), .Y(n3722) );
  CLKBUFX3 U2427 ( .A(n3786), .Y(n3723) );
  CLKBUFX3 U2428 ( .A(n3786), .Y(n3724) );
  CLKBUFX3 U2429 ( .A(n3786), .Y(n3725) );
  CLKBUFX3 U2430 ( .A(n3785), .Y(n3726) );
  CLKBUFX3 U2431 ( .A(n3785), .Y(n3727) );
  CLKBUFX3 U2432 ( .A(n3785), .Y(n3728) );
  CLKBUFX3 U2433 ( .A(n3785), .Y(n3729) );
  CLKBUFX3 U2434 ( .A(n3800), .Y(n3730) );
  CLKBUFX3 U2435 ( .A(n3800), .Y(n3731) );
  CLKBUFX3 U2436 ( .A(n3789), .Y(n3732) );
  CLKBUFX3 U2437 ( .A(n3788), .Y(n3733) );
  CLKBUFX3 U2438 ( .A(n3801), .Y(n3734) );
  CLKBUFX3 U2439 ( .A(n3794), .Y(n3735) );
  CLKBUFX3 U2440 ( .A(n3793), .Y(n3736) );
  CLKBUFX3 U2441 ( .A(n3792), .Y(n3737) );
  CLKBUFX3 U2442 ( .A(n3801), .Y(n3738) );
  CLKBUFX3 U2443 ( .A(n3781), .Y(n3739) );
  CLKBUFX3 U2444 ( .A(n3796), .Y(n3740) );
  CLKBUFX3 U2445 ( .A(n3795), .Y(n3741) );
  CLKBUFX3 U2446 ( .A(n3784), .Y(n3742) );
  CLKBUFX3 U2447 ( .A(n3784), .Y(n3743) );
  CLKBUFX3 U2448 ( .A(n3784), .Y(n3744) );
  CLKBUFX3 U2449 ( .A(n3784), .Y(n3745) );
  CLKBUFX3 U2450 ( .A(n3801), .Y(n3746) );
  CLKBUFX3 U2451 ( .A(n3801), .Y(n3747) );
  CLKBUFX3 U2452 ( .A(n3791), .Y(n3748) );
  CLKBUFX3 U2453 ( .A(n3790), .Y(n3749) );
  CLKBUFX3 U2454 ( .A(n3802), .Y(n3750) );
  CLKBUFX3 U2455 ( .A(n3802), .Y(n3751) );
  CLKBUFX3 U2456 ( .A(n3670), .Y(n3752) );
  CLKBUFX3 U2457 ( .A(n3799), .Y(n3753) );
  CLKBUFX3 U2458 ( .A(n3802), .Y(n3754) );
  CLKBUFX3 U2459 ( .A(n3782), .Y(n3755) );
  CLKBUFX3 U2460 ( .A(n3784), .Y(n3756) );
  CLKBUFX3 U2461 ( .A(n4120), .Y(n3757) );
  CLKBUFX3 U2462 ( .A(n4120), .Y(n3758) );
  CLKBUFX3 U2463 ( .A(n3802), .Y(n3759) );
  CLKBUFX3 U2464 ( .A(n3803), .Y(n3760) );
  CLKBUFX3 U2465 ( .A(n3803), .Y(n3761) );
  CLKBUFX3 U2466 ( .A(n3669), .Y(n3762) );
  CLKBUFX3 U2467 ( .A(n3783), .Y(n3763) );
  CLKBUFX3 U2468 ( .A(n3783), .Y(n3764) );
  CLKBUFX3 U2469 ( .A(n3783), .Y(n3765) );
  CLKBUFX3 U2470 ( .A(n3782), .Y(n3766) );
  CLKBUFX3 U2471 ( .A(n3782), .Y(n3767) );
  CLKBUFX3 U2472 ( .A(n3782), .Y(n3768) );
  CLKBUFX3 U2473 ( .A(n3782), .Y(n3769) );
  CLKBUFX3 U2474 ( .A(n3804), .Y(n3770) );
  CLKBUFX3 U2475 ( .A(n3804), .Y(n3771) );
  CLKBUFX3 U2476 ( .A(n3803), .Y(n3772) );
  CLKBUFX3 U2477 ( .A(n3783), .Y(n3773) );
  CLKBUFX3 U2478 ( .A(n3781), .Y(n3774) );
  CLKBUFX3 U2479 ( .A(n3781), .Y(n3775) );
  CLKBUFX3 U2480 ( .A(n3781), .Y(n3776) );
  CLKBUFX3 U2481 ( .A(n3781), .Y(n3777) );
  CLKBUFX3 U2482 ( .A(n3804), .Y(n3778) );
  CLKBUFX3 U2483 ( .A(n3804), .Y(n3779) );
  CLKBUFX3 U2484 ( .A(n3783), .Y(n3780) );
  CLKBUFX3 U2485 ( .A(n3797), .Y(n3671) );
  CLKBUFX3 U2486 ( .A(n3802), .Y(n3672) );
  CLKBUFX3 U2487 ( .A(n4120), .Y(n3673) );
  CLKBUFX3 U2488 ( .A(n3623), .Y(n3597) );
  CLKBUFX3 U2489 ( .A(n3623), .Y(n3596) );
  CLKBUFX3 U2490 ( .A(n3624), .Y(n3629) );
  CLKBUFX3 U2491 ( .A(n3655), .Y(n3624) );
  CLKBUFX3 U2492 ( .A(N43), .Y(n3655) );
  INVX3 U2493 ( .A(n3809), .Y(n3807) );
  CLKBUFX3 U2494 ( .A(n4122), .Y(n3805) );
  CLKBUFX3 U2495 ( .A(n4112), .Y(n4113) );
  CLKBUFX3 U2496 ( .A(n4122), .Y(n3806) );
  CLKBUFX3 U2497 ( .A(n267), .Y(n3997) );
  CLKBUFX3 U2498 ( .A(n3960), .Y(n3992) );
  CLKBUFX3 U2499 ( .A(n3960), .Y(n3993) );
  CLKBUFX3 U2500 ( .A(n3960), .Y(n3994) );
  CLKBUFX3 U2501 ( .A(n3960), .Y(n3995) );
  CLKBUFX3 U2502 ( .A(n3960), .Y(n3996) );
  CLKBUFX3 U2503 ( .A(n3857), .Y(n3856) );
  CLKBUFX3 U2504 ( .A(n3870), .Y(n3869) );
  CLKBUFX3 U2505 ( .A(n283), .Y(n3882) );
  CLKBUFX3 U2506 ( .A(n3896), .Y(n3895) );
  CLKBUFX3 U2507 ( .A(n3909), .Y(n3908) );
  CLKBUFX3 U2508 ( .A(n3922), .Y(n3921) );
  CLKBUFX3 U2509 ( .A(n3935), .Y(n3934) );
  CLKBUFX3 U2510 ( .A(n3948), .Y(n3947) );
  INVX3 U2511 ( .A(n3235), .Y(n3808) );
  CLKBUFX3 U2512 ( .A(n3797), .Y(n3796) );
  CLKBUFX3 U2513 ( .A(n3797), .Y(n3795) );
  CLKBUFX3 U2514 ( .A(n3798), .Y(n3794) );
  CLKBUFX3 U2515 ( .A(n3798), .Y(n3793) );
  CLKBUFX3 U2516 ( .A(n3798), .Y(n3792) );
  CLKBUFX3 U2517 ( .A(n3799), .Y(n3791) );
  CLKBUFX3 U2518 ( .A(n3799), .Y(n3790) );
  CLKBUFX3 U2519 ( .A(n3799), .Y(n3789) );
  CLKBUFX3 U2520 ( .A(n3799), .Y(n3788) );
  CLKBUFX3 U2521 ( .A(n3800), .Y(n3787) );
  CLKBUFX3 U2522 ( .A(n3800), .Y(n3786) );
  CLKBUFX3 U2523 ( .A(n3800), .Y(n3785) );
  CLKBUFX3 U2524 ( .A(n3801), .Y(n3784) );
  CLKBUFX3 U2525 ( .A(n3803), .Y(n3783) );
  CLKBUFX3 U2526 ( .A(n3803), .Y(n3782) );
  CLKBUFX3 U2527 ( .A(n3804), .Y(n3781) );
  CLKBUFX3 U2528 ( .A(n3268), .Y(n4112) );
  OA21XL U2529 ( .A0(n102), .A1(n190), .B0(n3860), .Y(n3278) );
  CLKINVX1 U2530 ( .A(n3278), .Y(n195) );
  OA21XL U2531 ( .A0(n102), .A1(n139), .B0(n3872), .Y(n3279) );
  CLKINVX1 U2532 ( .A(n3279), .Y(n185) );
  NAND2BX2 U2533 ( .AN(n3668), .B(n269), .Y(n306) );
  NAND2X1 U2534 ( .A(n3808), .B(n199), .Y(n269) );
  CLKBUFX3 U2535 ( .A(n197), .Y(n4004) );
  CLKBUFX3 U2536 ( .A(n197), .Y(n4005) );
  CLKBUFX3 U2537 ( .A(n197), .Y(n4003) );
  CLKBUFX3 U2538 ( .A(n3811), .Y(n3809) );
  CLKBUFX3 U2539 ( .A(n205), .Y(n3999) );
  CLKBUFX3 U2540 ( .A(n208), .Y(n3998) );
  CLKBUFX3 U2541 ( .A(n267), .Y(n3960) );
  CLKBUFX3 U2542 ( .A(n284), .Y(n3870) );
  CLKBUFX3 U2543 ( .A(n285), .Y(n3857) );
  CLKBUFX3 U2544 ( .A(n282), .Y(n3896) );
  CLKBUFX3 U2545 ( .A(n280), .Y(n3909) );
  CLKBUFX3 U2546 ( .A(n278), .Y(n3922) );
  CLKBUFX3 U2547 ( .A(n276), .Y(n3935) );
  CLKBUFX3 U2548 ( .A(n274), .Y(n3948) );
  CLKBUFX3 U2549 ( .A(n3809), .Y(n3810) );
  NAND3X2 U2550 ( .A(n4118), .B(n4116), .C(n4114), .Y(n305) );
  CLKBUFX3 U2551 ( .A(n3285), .Y(n3287) );
  CLKBUFX3 U2552 ( .A(n3285), .Y(n3286) );
  CLKINVX1 U2553 ( .A(n270), .Y(n4121) );
  INVX3 U2554 ( .A(n4002), .Y(n4001) );
  CLKBUFX3 U2555 ( .A(n3214), .Y(n4028) );
  CLKBUFX3 U2556 ( .A(n3215), .Y(n4030) );
  CLKBUFX3 U2557 ( .A(n3216), .Y(n4032) );
  CLKBUFX3 U2558 ( .A(n3205), .Y(n4034) );
  CLKBUFX3 U2559 ( .A(n3206), .Y(n4036) );
  CLKBUFX3 U2560 ( .A(n3207), .Y(n4038) );
  CLKBUFX3 U2561 ( .A(n3208), .Y(n4040) );
  CLKBUFX3 U2562 ( .A(n3217), .Y(n4044) );
  CLKBUFX3 U2563 ( .A(n3218), .Y(n4047) );
  CLKBUFX3 U2564 ( .A(n3203), .Y(n4049) );
  CLKBUFX3 U2565 ( .A(n3204), .Y(n4051) );
  CLKBUFX3 U2566 ( .A(n3210), .Y(n4053) );
  CLKBUFX3 U2567 ( .A(n3211), .Y(n4055) );
  CLKBUFX3 U2568 ( .A(n3212), .Y(n4057) );
  CLKBUFX3 U2569 ( .A(n3213), .Y(n4059) );
  CLKBUFX3 U2570 ( .A(n3219), .Y(n4062) );
  CLKBUFX3 U2571 ( .A(n3220), .Y(n4065) );
  CLKBUFX3 U2572 ( .A(n3221), .Y(n4068) );
  CLKBUFX3 U2573 ( .A(n3222), .Y(n4071) );
  CLKBUFX3 U2574 ( .A(n3223), .Y(n4074) );
  CLKBUFX3 U2575 ( .A(n3224), .Y(n4077) );
  CLKBUFX3 U2576 ( .A(n3225), .Y(n4080) );
  CLKBUFX3 U2577 ( .A(n3226), .Y(n4083) );
  CLKBUFX3 U2578 ( .A(n3227), .Y(n4086) );
  CLKBUFX3 U2579 ( .A(n3228), .Y(n4089) );
  CLKBUFX3 U2580 ( .A(n3229), .Y(n4092) );
  CLKBUFX3 U2581 ( .A(n3230), .Y(n4095) );
  CLKBUFX3 U2582 ( .A(n3231), .Y(n4098) );
  CLKBUFX3 U2583 ( .A(n3232), .Y(n4101) );
  CLKBUFX3 U2584 ( .A(n3233), .Y(n4104) );
  CLKBUFX3 U2585 ( .A(n3234), .Y(n4107) );
  CLKBUFX3 U2586 ( .A(n3217), .Y(n4045) );
  CLKBUFX3 U2587 ( .A(n3218), .Y(n4048) );
  CLKBUFX3 U2588 ( .A(n3203), .Y(n4050) );
  CLKBUFX3 U2589 ( .A(n3204), .Y(n4052) );
  CLKBUFX3 U2590 ( .A(n3210), .Y(n4054) );
  CLKBUFX3 U2591 ( .A(n3211), .Y(n4056) );
  CLKBUFX3 U2592 ( .A(n3212), .Y(n4058) );
  CLKBUFX3 U2593 ( .A(n3213), .Y(n4060) );
  CLKBUFX3 U2594 ( .A(n3219), .Y(n4063) );
  CLKBUFX3 U2595 ( .A(n3220), .Y(n4066) );
  CLKBUFX3 U2596 ( .A(n3221), .Y(n4069) );
  CLKBUFX3 U2597 ( .A(n3222), .Y(n4072) );
  CLKBUFX3 U2598 ( .A(n3223), .Y(n4075) );
  CLKBUFX3 U2599 ( .A(n3224), .Y(n4078) );
  CLKBUFX3 U2600 ( .A(n3225), .Y(n4081) );
  CLKBUFX3 U2601 ( .A(n3226), .Y(n4084) );
  CLKBUFX3 U2602 ( .A(n3227), .Y(n4087) );
  CLKBUFX3 U2603 ( .A(n3228), .Y(n4090) );
  CLKBUFX3 U2604 ( .A(n3229), .Y(n4093) );
  CLKBUFX3 U2605 ( .A(n3230), .Y(n4096) );
  CLKBUFX3 U2606 ( .A(n3231), .Y(n4099) );
  CLKBUFX3 U2607 ( .A(n3232), .Y(n4102) );
  CLKBUFX3 U2608 ( .A(n3233), .Y(n4105) );
  CLKBUFX3 U2609 ( .A(n3234), .Y(n4108) );
  CLKBUFX3 U2610 ( .A(n3214), .Y(n4029) );
  CLKBUFX3 U2611 ( .A(n3215), .Y(n4031) );
  CLKBUFX3 U2612 ( .A(n3216), .Y(n4033) );
  CLKBUFX3 U2613 ( .A(n3205), .Y(n4035) );
  CLKBUFX3 U2614 ( .A(n3206), .Y(n4037) );
  CLKBUFX3 U2615 ( .A(n3207), .Y(n4039) );
  CLKBUFX3 U2616 ( .A(n3208), .Y(n4041) );
  CLKBUFX3 U2617 ( .A(N46), .Y(n3289) );
  CLKBUFX3 U2618 ( .A(N46), .Y(n3288) );
  CLKBUFX3 U2619 ( .A(n3209), .Y(n4111) );
  CLKBUFX3 U2620 ( .A(n3209), .Y(n4110) );
  CLKBUFX3 U2621 ( .A(n3669), .Y(n3797) );
  CLKBUFX3 U2622 ( .A(n3669), .Y(n3798) );
  CLKBUFX3 U2623 ( .A(n4120), .Y(n3799) );
  CLKBUFX3 U2624 ( .A(n3670), .Y(n3800) );
  CLKBUFX3 U2625 ( .A(n3670), .Y(n3801) );
  CLKBUFX3 U2626 ( .A(n3670), .Y(n3802) );
  CLKBUFX3 U2627 ( .A(n3670), .Y(n3803) );
  CLKBUFX3 U2628 ( .A(n3669), .Y(n3804) );
  NOR4X1 U2629 ( .A(n394), .B(n395), .C(n396), .D(n397), .Y(n368) );
  NOR4X1 U2630 ( .A(n386), .B(n387), .C(n388), .D(n389), .Y(n369) );
  XNOR2X1 U2631 ( .A(n4127), .B(N210), .Y(n375) );
  XNOR2X1 U2632 ( .A(n4143), .B(N226), .Y(n389) );
  XNOR2X1 U2633 ( .A(n4142), .B(N225), .Y(n397) );
  XNOR2X1 U2634 ( .A(n4126), .B(N209), .Y(n374) );
  XNOR2X1 U2635 ( .A(n4124), .B(N207), .Y(n388) );
  XNOR2X1 U2636 ( .A(n4146), .B(N229), .Y(n396) );
  XNOR2X1 U2637 ( .A(n4125), .B(N208), .Y(n373) );
  XNOR2X1 U2638 ( .A(n4130), .B(N213), .Y(n387) );
  XNOR2X1 U2639 ( .A(n4144), .B(N227), .Y(n395) );
  NOR4X1 U2640 ( .A(n379), .B(n380), .C(n381), .D(n382), .Y(n370) );
  XNOR2X1 U2641 ( .A(n4132), .B(N215), .Y(n380) );
  NAND3X1 U2642 ( .A(n383), .B(n384), .C(n385), .Y(n379) );
  XNOR2X1 U2643 ( .A(n4141), .B(N224), .Y(n381) );
  AOI21X1 U2644 ( .A0(n265), .A1(n199), .B0(n260), .Y(n261) );
  NAND3X2 U2645 ( .A(n4119), .B(n4115), .C(n4116), .Y(n101) );
  OAI21X1 U2646 ( .A0(n4123), .A1(n200), .B0(n4000), .Y(n202) );
  CLKINVX1 U2647 ( .A(n199), .Y(n4123) );
  NAND2X1 U2648 ( .A(N233), .B(n258), .Y(n208) );
  AOI211X1 U2649 ( .A0(n291), .A1(n292), .B0(n4304), .C0(n289), .Y(n3171) );
  NOR2X1 U2650 ( .A(n260), .B(n288), .Y(n291) );
  OAI21XL U2651 ( .A0(n4172), .A1(n269), .B0(n290), .Y(n292) );
  NOR2X1 U2652 ( .A(n139), .B(n3667), .Y(n284) );
  NOR2X1 U2653 ( .A(n190), .B(n3667), .Y(n285) );
  NOR2X1 U2654 ( .A(n315), .B(n3667), .Y(n282) );
  NOR2X1 U2655 ( .A(n313), .B(n3667), .Y(n280) );
  NOR2X1 U2656 ( .A(n311), .B(n3667), .Y(n278) );
  NOR2X1 U2657 ( .A(n309), .B(n3667), .Y(n276) );
  NOR2X1 U2658 ( .A(n305), .B(n3667), .Y(n274) );
  NOR2X1 U2659 ( .A(n3667), .B(n101), .Y(n283) );
  NOR2X1 U2660 ( .A(n261), .B(n260), .Y(n258) );
  CLKBUFX3 U2661 ( .A(n308), .Y(n3668) );
  CLKINVX1 U2662 ( .A(n1713), .Y(n3811) );
  NAND3X2 U2663 ( .A(n4116), .B(n4115), .C(n4118), .Y(n315) );
  NAND3X2 U2664 ( .A(n4119), .B(n4117), .C(n4114), .Y(n313) );
  NAND3X2 U2665 ( .A(n4118), .B(n4117), .C(n4114), .Y(n311) );
  NAND3X2 U2666 ( .A(n4116), .B(n4119), .C(n4114), .Y(n309) );
  CLKINVX1 U2667 ( .A(N233), .Y(n4172) );
  CLKINVX1 U2668 ( .A(n260), .Y(n4303) );
  NAND3X1 U2669 ( .A(n4303), .B(n3667), .C(n295), .Y(n270) );
  NAND2X1 U2670 ( .A(n4000), .B(n200), .Y(n265) );
  AND3X2 U2671 ( .A(n4305), .B(n290), .C(n295), .Y(n289) );
  CLKINVX1 U2672 ( .A(n288), .Y(n4305) );
  CLKBUFX3 U2673 ( .A(n3281), .Y(n4002) );
  CLKINVX1 U2674 ( .A(n3667), .Y(n4304) );
  CLKBUFX3 U2675 ( .A(n3217), .Y(n4043) );
  CLKBUFX3 U2676 ( .A(n3218), .Y(n4046) );
  CLKBUFX3 U2677 ( .A(n3219), .Y(n4061) );
  CLKBUFX3 U2678 ( .A(n3220), .Y(n4064) );
  CLKBUFX3 U2679 ( .A(n3221), .Y(n4067) );
  CLKBUFX3 U2680 ( .A(n3222), .Y(n4070) );
  CLKBUFX3 U2681 ( .A(n3223), .Y(n4073) );
  CLKBUFX3 U2682 ( .A(n3224), .Y(n4076) );
  CLKBUFX3 U2683 ( .A(n3225), .Y(n4079) );
  CLKBUFX3 U2684 ( .A(n3226), .Y(n4082) );
  CLKBUFX3 U2685 ( .A(n3227), .Y(n4085) );
  CLKBUFX3 U2686 ( .A(n3228), .Y(n4088) );
  CLKBUFX3 U2687 ( .A(n3229), .Y(n4091) );
  CLKBUFX3 U2688 ( .A(n3230), .Y(n4094) );
  CLKBUFX3 U2689 ( .A(n3231), .Y(n4097) );
  CLKBUFX3 U2690 ( .A(n3232), .Y(n4100) );
  CLKBUFX3 U2691 ( .A(n3233), .Y(n4103) );
  CLKBUFX3 U2692 ( .A(n3234), .Y(n4106) );
  OAI2BB1X1 U2693 ( .A0N(n3810), .A1N(n198), .B0(n3667), .Y(n3172) );
  CLKBUFX3 U2694 ( .A(n3238), .Y(n3669) );
  CLKBUFX3 U2695 ( .A(n3237), .Y(n3670) );
  OAI222XL U2696 ( .A0(n402), .A1(n4113), .B0(n4109), .B1(n4030), .C0(n3884), 
        .C1(n4244), .Y(n2433) );
  OAI222XL U2697 ( .A0(n404), .A1(n4113), .B0(n4109), .B1(n4034), .C0(n3884), 
        .C1(n4242), .Y(n2431) );
  OAI222XL U2698 ( .A0(n405), .A1(n4113), .B0(n4109), .B1(n4036), .C0(n3885), 
        .C1(n4241), .Y(n2430) );
  OAI222XL U2699 ( .A0(n407), .A1(n4112), .B0(n4109), .B1(n4040), .C0(n3885), 
        .C1(n4239), .Y(n2428) );
  OAI222XL U2700 ( .A0(n1671), .A1(n4112), .B0(n4109), .B1(n4044), .C0(n3890), 
        .C1(n4270), .Y(n2459) );
  OAI222XL U2701 ( .A0(n1672), .A1(n4112), .B0(n4109), .B1(n4047), .C0(n3890), 
        .C1(n4269), .Y(n2458) );
  OAI222XL U2702 ( .A0(n1673), .A1(n4112), .B0(n4109), .B1(n4049), .C0(n3890), 
        .C1(n4268), .Y(n2457) );
  OAI222XL U2703 ( .A0(n1674), .A1(n4112), .B0(n4109), .B1(n4051), .C0(n3890), 
        .C1(n4267), .Y(n2456) );
  OAI222XL U2704 ( .A0(n1675), .A1(n4112), .B0(n4109), .B1(n4053), .C0(n3890), 
        .C1(n4266), .Y(n2455) );
  OAI222XL U2705 ( .A0(n1676), .A1(n4112), .B0(n4109), .B1(n4055), .C0(n3890), 
        .C1(n4265), .Y(n2454) );
  OAI222XL U2706 ( .A0(n1677), .A1(n4112), .B0(n4109), .B1(n4057), .C0(n3890), 
        .C1(n4264), .Y(n2453) );
  OAI222XL U2707 ( .A0(n1678), .A1(n4113), .B0(n4109), .B1(n4059), .C0(n3890), 
        .C1(n4263), .Y(n2452) );
  OAI222XL U2708 ( .A0(n1679), .A1(n4113), .B0(n4109), .B1(n4062), .C0(n3890), 
        .C1(n4262), .Y(n2451) );
  OAI222XL U2709 ( .A0(n1680), .A1(n4113), .B0(n4109), .B1(n4065), .C0(n3890), 
        .C1(n4261), .Y(n2450) );
  OAI222XL U2710 ( .A0(n1681), .A1(n4113), .B0(n4109), .B1(n4068), .C0(n3890), 
        .C1(n4260), .Y(n2449) );
  OAI222XL U2711 ( .A0(n1682), .A1(n4113), .B0(n4109), .B1(n4071), .C0(n3890), 
        .C1(n4259), .Y(n2448) );
  OAI222XL U2712 ( .A0(n1683), .A1(n4113), .B0(n4109), .B1(n4074), .C0(n3891), 
        .C1(n4258), .Y(n2447) );
  OAI222XL U2713 ( .A0(n1684), .A1(n4113), .B0(n4109), .B1(n4077), .C0(n3891), 
        .C1(n4257), .Y(n2446) );
  OAI222XL U2714 ( .A0(n1685), .A1(n4113), .B0(n4109), .B1(n4080), .C0(n3891), 
        .C1(n4256), .Y(n2445) );
  OAI222XL U2715 ( .A0(n1686), .A1(n4113), .B0(n4109), .B1(n4083), .C0(n3891), 
        .C1(n4255), .Y(n2444) );
  OAI222XL U2716 ( .A0(n1687), .A1(n4113), .B0(n4109), .B1(n4086), .C0(n3891), 
        .C1(n4254), .Y(n2443) );
  OAI222XL U2717 ( .A0(n1688), .A1(n4113), .B0(n4109), .B1(n4089), .C0(n3891), 
        .C1(n4253), .Y(n2442) );
  OAI222XL U2718 ( .A0(n1689), .A1(n4113), .B0(n4109), .B1(n4092), .C0(n3891), 
        .C1(n4252), .Y(n2441) );
  OAI222XL U2719 ( .A0(n1690), .A1(n4113), .B0(n4109), .B1(n4095), .C0(n3891), 
        .C1(n4251), .Y(n2440) );
  OAI222XL U2720 ( .A0(n1691), .A1(n4113), .B0(n4109), .B1(n4098), .C0(n3891), 
        .C1(n4250), .Y(n2439) );
  OAI222XL U2721 ( .A0(n1692), .A1(n4113), .B0(n4109), .B1(n4101), .C0(n3891), 
        .C1(n4249), .Y(n2438) );
  OAI222XL U2722 ( .A0(n1693), .A1(n4113), .B0(n4109), .B1(n4104), .C0(n3891), 
        .C1(n4248), .Y(n2437) );
  OAI222XL U2723 ( .A0(n1694), .A1(n4113), .B0(n4109), .B1(n4107), .C0(n3891), 
        .C1(n4247), .Y(n2436) );
  OAI222XL U2724 ( .A0(n1695), .A1(n4113), .B0(n4110), .B1(n4109), .C0(n3884), 
        .C1(n4246), .Y(n2435) );
  OAI222XL U2725 ( .A0(n504), .A1(n3175), .B0(n4043), .B1(n3819), .C0(n4270), 
        .C1(n3902), .Y(n2331) );
  OAI222XL U2726 ( .A0(n505), .A1(n3175), .B0(n4046), .B1(n3818), .C0(n4269), 
        .C1(n3900), .Y(n2330) );
  OAI222XL U2727 ( .A0(n506), .A1(n3175), .B0(n3203), .B1(n359), .C0(n4268), 
        .C1(n3904), .Y(n2329) );
  OAI222XL U2728 ( .A0(n507), .A1(n3175), .B0(n3204), .B1(n359), .C0(n4267), 
        .C1(n3900), .Y(n2328) );
  OAI222XL U2729 ( .A0(n508), .A1(n3175), .B0(n3210), .B1(n359), .C0(n4266), 
        .C1(n3901), .Y(n2327) );
  OAI222XL U2730 ( .A0(n509), .A1(n3175), .B0(n3211), .B1(n359), .C0(n4265), 
        .C1(n3900), .Y(n2326) );
  OAI222XL U2731 ( .A0(n510), .A1(n3175), .B0(n3212), .B1(n359), .C0(n4264), 
        .C1(n3900), .Y(n2325) );
  OAI222XL U2732 ( .A0(n511), .A1(n3175), .B0(n3213), .B1(n359), .C0(n4263), 
        .C1(n3900), .Y(n2324) );
  OAI222XL U2733 ( .A0(n512), .A1(n3175), .B0(n4061), .B1(n3819), .C0(n4262), 
        .C1(n3900), .Y(n2323) );
  OAI222XL U2734 ( .A0(n513), .A1(n3175), .B0(n4064), .B1(n3819), .C0(n4261), 
        .C1(n3900), .Y(n2322) );
  OAI222XL U2735 ( .A0(n514), .A1(n3175), .B0(n4067), .B1(n3819), .C0(n4260), 
        .C1(n3900), .Y(n2321) );
  OAI222XL U2736 ( .A0(n515), .A1(n3175), .B0(n4070), .B1(n3819), .C0(n4259), 
        .C1(n3900), .Y(n2320) );
  OAI222XL U2737 ( .A0(n516), .A1(n3175), .B0(n4073), .B1(n3819), .C0(n4258), 
        .C1(n3900), .Y(n2319) );
  OAI222XL U2738 ( .A0(n517), .A1(n3175), .B0(n4076), .B1(n3819), .C0(n4257), 
        .C1(n3900), .Y(n2318) );
  OAI222XL U2739 ( .A0(n518), .A1(n3175), .B0(n4079), .B1(n3819), .C0(n4256), 
        .C1(n3900), .Y(n2317) );
  OAI222XL U2740 ( .A0(n519), .A1(n3175), .B0(n4082), .B1(n3819), .C0(n4255), 
        .C1(n3900), .Y(n2316) );
  OAI222XL U2741 ( .A0(n520), .A1(n3175), .B0(n4085), .B1(n3819), .C0(n4254), 
        .C1(n3900), .Y(n2315) );
  OAI222XL U2742 ( .A0(n521), .A1(n3175), .B0(n4088), .B1(n3819), .C0(n4253), 
        .C1(n3900), .Y(n2314) );
  OAI222XL U2743 ( .A0(n522), .A1(n3175), .B0(n4091), .B1(n3819), .C0(n4252), 
        .C1(n3900), .Y(n2313) );
  OAI222XL U2744 ( .A0(n523), .A1(n3175), .B0(n4094), .B1(n3819), .C0(n4251), 
        .C1(n3901), .Y(n2312) );
  OAI222XL U2745 ( .A0(n524), .A1(n3175), .B0(n4097), .B1(n3818), .C0(n4250), 
        .C1(n3900), .Y(n2311) );
  OAI222XL U2746 ( .A0(n525), .A1(n3175), .B0(n4100), .B1(n3818), .C0(n4249), 
        .C1(n3901), .Y(n2310) );
  OAI222XL U2747 ( .A0(n526), .A1(n3175), .B0(n4103), .B1(n3818), .C0(n4248), 
        .C1(n3901), .Y(n2309) );
  OAI222XL U2748 ( .A0(n527), .A1(n3175), .B0(n4106), .B1(n3818), .C0(n4247), 
        .C1(n3901), .Y(n2308) );
  OAI222XL U2749 ( .A0(n528), .A1(n3175), .B0(n4111), .B1(n3818), .C0(n4246), 
        .C1(n3901), .Y(n2307) );
  OAI222XL U2750 ( .A0(n529), .A1(n3175), .B0(n4028), .B1(n3818), .C0(n4245), 
        .C1(n3901), .Y(n2306) );
  OAI222XL U2751 ( .A0(n530), .A1(n3175), .B0(n4030), .B1(n3818), .C0(n4244), 
        .C1(n3901), .Y(n2305) );
  OAI222XL U2752 ( .A0(n531), .A1(n3175), .B0(n4032), .B1(n3818), .C0(n4243), 
        .C1(n3901), .Y(n2304) );
  OAI222XL U2753 ( .A0(n532), .A1(n3175), .B0(n4034), .B1(n3818), .C0(n4242), 
        .C1(n3901), .Y(n2303) );
  OAI222XL U2754 ( .A0(n533), .A1(n3175), .B0(n4036), .B1(n3818), .C0(n4241), 
        .C1(n3901), .Y(n2302) );
  OAI222XL U2755 ( .A0(n534), .A1(n3175), .B0(n4038), .B1(n3818), .C0(n4240), 
        .C1(n3901), .Y(n2301) );
  OAI222XL U2756 ( .A0(n535), .A1(n3175), .B0(n4040), .B1(n3818), .C0(n4239), 
        .C1(n3901), .Y(n2300) );
  OAI222XL U2757 ( .A0(n632), .A1(n3183), .B0(n4045), .B1(n3827), .C0(n4270), 
        .C1(n3912), .Y(n2203) );
  OAI222XL U2758 ( .A0(n633), .A1(n3183), .B0(n4048), .B1(n3826), .C0(n4269), 
        .C1(n3913), .Y(n2202) );
  OAI222XL U2759 ( .A0(n634), .A1(n3183), .B0(n4050), .B1(n351), .C0(n4268), 
        .C1(n3910), .Y(n2201) );
  OAI222XL U2760 ( .A0(n635), .A1(n3183), .B0(n4052), .B1(n351), .C0(n4267), 
        .C1(n3910), .Y(n2200) );
  OAI222XL U2761 ( .A0(n636), .A1(n3183), .B0(n4054), .B1(n351), .C0(n4266), 
        .C1(n3914), .Y(n2199) );
  OAI222XL U2762 ( .A0(n637), .A1(n3183), .B0(n4056), .B1(n351), .C0(n4265), 
        .C1(n3913), .Y(n2198) );
  OAI222XL U2763 ( .A0(n638), .A1(n3183), .B0(n4058), .B1(n351), .C0(n4264), 
        .C1(n3913), .Y(n2197) );
  OAI222XL U2764 ( .A0(n639), .A1(n3183), .B0(n4060), .B1(n351), .C0(n4263), 
        .C1(n3913), .Y(n2196) );
  OAI222XL U2765 ( .A0(n640), .A1(n3183), .B0(n4063), .B1(n3827), .C0(n4262), 
        .C1(n3913), .Y(n2195) );
  OAI222XL U2766 ( .A0(n641), .A1(n3183), .B0(n4066), .B1(n3827), .C0(n4261), 
        .C1(n3913), .Y(n2194) );
  OAI222XL U2767 ( .A0(n642), .A1(n3183), .B0(n4069), .B1(n3827), .C0(n4260), 
        .C1(n3913), .Y(n2193) );
  OAI222XL U2768 ( .A0(n643), .A1(n3183), .B0(n4072), .B1(n3827), .C0(n4259), 
        .C1(n3913), .Y(n2192) );
  OAI222XL U2769 ( .A0(n644), .A1(n3183), .B0(n4075), .B1(n3827), .C0(n4258), 
        .C1(n3913), .Y(n2191) );
  OAI222XL U2770 ( .A0(n645), .A1(n3183), .B0(n4078), .B1(n3827), .C0(n4257), 
        .C1(n3913), .Y(n2190) );
  OAI222XL U2771 ( .A0(n646), .A1(n3183), .B0(n4081), .B1(n3827), .C0(n4256), 
        .C1(n3913), .Y(n2189) );
  OAI222XL U2772 ( .A0(n647), .A1(n3183), .B0(n4084), .B1(n3827), .C0(n4255), 
        .C1(n3913), .Y(n2188) );
  OAI222XL U2773 ( .A0(n648), .A1(n3183), .B0(n4087), .B1(n3827), .C0(n4254), 
        .C1(n3913), .Y(n2187) );
  OAI222XL U2774 ( .A0(n649), .A1(n3183), .B0(n4090), .B1(n3827), .C0(n4253), 
        .C1(n3913), .Y(n2186) );
  OAI222XL U2775 ( .A0(n650), .A1(n3183), .B0(n4093), .B1(n3827), .C0(n4252), 
        .C1(n3913), .Y(n2185) );
  OAI222XL U2776 ( .A0(n651), .A1(n3183), .B0(n4096), .B1(n3827), .C0(n4251), 
        .C1(n3914), .Y(n2184) );
  OAI222XL U2777 ( .A0(n652), .A1(n3183), .B0(n4099), .B1(n3826), .C0(n4250), 
        .C1(n3913), .Y(n2183) );
  OAI222XL U2778 ( .A0(n653), .A1(n3183), .B0(n4102), .B1(n3826), .C0(n4249), 
        .C1(n3914), .Y(n2182) );
  OAI222XL U2779 ( .A0(n654), .A1(n3183), .B0(n4105), .B1(n3826), .C0(n4248), 
        .C1(n3914), .Y(n2181) );
  OAI222XL U2780 ( .A0(n655), .A1(n3183), .B0(n4108), .B1(n3826), .C0(n4247), 
        .C1(n3914), .Y(n2180) );
  OAI222XL U2781 ( .A0(n656), .A1(n3183), .B0(n4110), .B1(n3826), .C0(n4246), 
        .C1(n3914), .Y(n2179) );
  OAI222XL U2782 ( .A0(n657), .A1(n3183), .B0(n4029), .B1(n3826), .C0(n4245), 
        .C1(n3914), .Y(n2178) );
  OAI222XL U2783 ( .A0(n658), .A1(n3183), .B0(n4031), .B1(n3826), .C0(n4244), 
        .C1(n3914), .Y(n2177) );
  OAI222XL U2784 ( .A0(n659), .A1(n3183), .B0(n4033), .B1(n3826), .C0(n4243), 
        .C1(n3914), .Y(n2176) );
  OAI222XL U2785 ( .A0(n660), .A1(n3183), .B0(n4035), .B1(n3826), .C0(n4242), 
        .C1(n3914), .Y(n2175) );
  OAI222XL U2786 ( .A0(n661), .A1(n3183), .B0(n4037), .B1(n3826), .C0(n4241), 
        .C1(n3914), .Y(n2174) );
  OAI222XL U2787 ( .A0(n662), .A1(n3183), .B0(n4039), .B1(n3826), .C0(n4240), 
        .C1(n3914), .Y(n2173) );
  OAI222XL U2788 ( .A0(n663), .A1(n3183), .B0(n4041), .B1(n3826), .C0(n4239), 
        .C1(n3914), .Y(n2172) );
  OAI222XL U2789 ( .A0(n760), .A1(n3181), .B0(n4045), .B1(n3835), .C0(n4270), 
        .C1(n3925), .Y(n2075) );
  OAI222XL U2790 ( .A0(n761), .A1(n3181), .B0(n4048), .B1(n3834), .C0(n4269), 
        .C1(n3926), .Y(n2074) );
  OAI222XL U2791 ( .A0(n762), .A1(n3181), .B0(n4050), .B1(n343), .C0(n4268), 
        .C1(n3923), .Y(n2073) );
  OAI222XL U2792 ( .A0(n763), .A1(n3181), .B0(n4052), .B1(n343), .C0(n4267), 
        .C1(n3923), .Y(n2072) );
  OAI222XL U2793 ( .A0(n764), .A1(n3181), .B0(n4054), .B1(n343), .C0(n4266), 
        .C1(n3927), .Y(n2071) );
  OAI222XL U2794 ( .A0(n765), .A1(n3181), .B0(n4056), .B1(n343), .C0(n4265), 
        .C1(n3926), .Y(n2070) );
  OAI222XL U2795 ( .A0(n766), .A1(n3181), .B0(n4058), .B1(n343), .C0(n4264), 
        .C1(n3926), .Y(n2069) );
  OAI222XL U2796 ( .A0(n767), .A1(n3181), .B0(n4060), .B1(n343), .C0(n4263), 
        .C1(n3926), .Y(n2068) );
  OAI222XL U2797 ( .A0(n768), .A1(n3181), .B0(n4063), .B1(n3835), .C0(n4262), 
        .C1(n3926), .Y(n2067) );
  OAI222XL U2798 ( .A0(n769), .A1(n3181), .B0(n4066), .B1(n3835), .C0(n4261), 
        .C1(n3926), .Y(n2066) );
  OAI222XL U2799 ( .A0(n770), .A1(n3181), .B0(n4069), .B1(n3835), .C0(n4260), 
        .C1(n3926), .Y(n2065) );
  OAI222XL U2800 ( .A0(n771), .A1(n3181), .B0(n4072), .B1(n3835), .C0(n4259), 
        .C1(n3926), .Y(n2064) );
  OAI222XL U2801 ( .A0(n772), .A1(n3181), .B0(n4075), .B1(n3835), .C0(n4258), 
        .C1(n3926), .Y(n2063) );
  OAI222XL U2802 ( .A0(n773), .A1(n3181), .B0(n4078), .B1(n3835), .C0(n4257), 
        .C1(n3926), .Y(n2062) );
  OAI222XL U2803 ( .A0(n774), .A1(n3181), .B0(n4081), .B1(n3835), .C0(n4256), 
        .C1(n3926), .Y(n2061) );
  OAI222XL U2804 ( .A0(n775), .A1(n3181), .B0(n4084), .B1(n3835), .C0(n4255), 
        .C1(n3926), .Y(n2060) );
  OAI222XL U2805 ( .A0(n776), .A1(n3181), .B0(n4087), .B1(n3835), .C0(n4254), 
        .C1(n3926), .Y(n2059) );
  OAI222XL U2806 ( .A0(n777), .A1(n3181), .B0(n4090), .B1(n3835), .C0(n4253), 
        .C1(n3926), .Y(n2058) );
  OAI222XL U2807 ( .A0(n778), .A1(n3181), .B0(n4093), .B1(n3835), .C0(n4252), 
        .C1(n3926), .Y(n2057) );
  OAI222XL U2808 ( .A0(n779), .A1(n3181), .B0(n4096), .B1(n3835), .C0(n4251), 
        .C1(n3927), .Y(n2056) );
  OAI222XL U2809 ( .A0(n780), .A1(n3181), .B0(n4099), .B1(n3834), .C0(n4250), 
        .C1(n3926), .Y(n2055) );
  OAI222XL U2810 ( .A0(n781), .A1(n3181), .B0(n4102), .B1(n3834), .C0(n4249), 
        .C1(n3927), .Y(n2054) );
  OAI222XL U2811 ( .A0(n782), .A1(n3181), .B0(n4105), .B1(n3834), .C0(n4248), 
        .C1(n3927), .Y(n2053) );
  OAI222XL U2812 ( .A0(n783), .A1(n3181), .B0(n4108), .B1(n3834), .C0(n4247), 
        .C1(n3927), .Y(n2052) );
  OAI222XL U2813 ( .A0(n784), .A1(n3181), .B0(n4111), .B1(n3834), .C0(n4246), 
        .C1(n3927), .Y(n2051) );
  OAI222XL U2814 ( .A0(n785), .A1(n3181), .B0(n4029), .B1(n3834), .C0(n4245), 
        .C1(n3927), .Y(n2050) );
  OAI222XL U2815 ( .A0(n786), .A1(n3181), .B0(n4031), .B1(n3834), .C0(n4244), 
        .C1(n3927), .Y(n2049) );
  OAI222XL U2816 ( .A0(n787), .A1(n3181), .B0(n4033), .B1(n3834), .C0(n4243), 
        .C1(n3927), .Y(n2048) );
  OAI222XL U2817 ( .A0(n788), .A1(n3181), .B0(n4035), .B1(n3834), .C0(n4242), 
        .C1(n3927), .Y(n2047) );
  OAI222XL U2818 ( .A0(n789), .A1(n3181), .B0(n4037), .B1(n3834), .C0(n4241), 
        .C1(n3927), .Y(n2046) );
  OAI222XL U2819 ( .A0(n790), .A1(n3181), .B0(n4039), .B1(n3834), .C0(n4240), 
        .C1(n3927), .Y(n2045) );
  OAI222XL U2820 ( .A0(n791), .A1(n3181), .B0(n4041), .B1(n3834), .C0(n4239), 
        .C1(n3927), .Y(n2044) );
  OAI222XL U2821 ( .A0(n888), .A1(n3179), .B0(n4045), .B1(n3843), .C0(n4270), 
        .C1(n3938), .Y(n1947) );
  OAI222XL U2822 ( .A0(n889), .A1(n3179), .B0(n4048), .B1(n3842), .C0(n4269), 
        .C1(n3939), .Y(n1946) );
  OAI222XL U2823 ( .A0(n890), .A1(n3179), .B0(n4050), .B1(n335), .C0(n4268), 
        .C1(n3942), .Y(n1945) );
  OAI222XL U2824 ( .A0(n891), .A1(n3179), .B0(n4052), .B1(n335), .C0(n4267), 
        .C1(n3936), .Y(n1944) );
  OAI222XL U2825 ( .A0(n892), .A1(n3179), .B0(n4054), .B1(n335), .C0(n4266), 
        .C1(n3940), .Y(n1943) );
  OAI222XL U2826 ( .A0(n893), .A1(n3179), .B0(n4056), .B1(n335), .C0(n4265), 
        .C1(n3939), .Y(n1942) );
  OAI222XL U2827 ( .A0(n894), .A1(n3179), .B0(n4058), .B1(n335), .C0(n4264), 
        .C1(n3939), .Y(n1941) );
  OAI222XL U2828 ( .A0(n895), .A1(n3179), .B0(n4060), .B1(n335), .C0(n4263), 
        .C1(n3939), .Y(n1940) );
  OAI222XL U2829 ( .A0(n896), .A1(n3179), .B0(n4063), .B1(n3843), .C0(n4262), 
        .C1(n3939), .Y(n1939) );
  OAI222XL U2830 ( .A0(n897), .A1(n3179), .B0(n4066), .B1(n3843), .C0(n4261), 
        .C1(n3939), .Y(n1938) );
  OAI222XL U2831 ( .A0(n898), .A1(n3179), .B0(n4069), .B1(n3843), .C0(n4260), 
        .C1(n3939), .Y(n1937) );
  OAI222XL U2832 ( .A0(n899), .A1(n3179), .B0(n4072), .B1(n3843), .C0(n4259), 
        .C1(n3939), .Y(n1936) );
  OAI222XL U2833 ( .A0(n900), .A1(n3179), .B0(n4075), .B1(n3843), .C0(n4258), 
        .C1(n3939), .Y(n1935) );
  OAI222XL U2834 ( .A0(n901), .A1(n3179), .B0(n4078), .B1(n3843), .C0(n4257), 
        .C1(n3939), .Y(n1934) );
  OAI222XL U2835 ( .A0(n902), .A1(n3179), .B0(n4081), .B1(n3843), .C0(n4256), 
        .C1(n3939), .Y(n1933) );
  OAI222XL U2836 ( .A0(n903), .A1(n3179), .B0(n4084), .B1(n3843), .C0(n4255), 
        .C1(n3939), .Y(n1932) );
  OAI222XL U2837 ( .A0(n904), .A1(n3179), .B0(n4087), .B1(n3843), .C0(n4254), 
        .C1(n3939), .Y(n1931) );
  OAI222XL U2838 ( .A0(n905), .A1(n3179), .B0(n4090), .B1(n3843), .C0(n4253), 
        .C1(n3939), .Y(n1930) );
  OAI222XL U2839 ( .A0(n906), .A1(n3179), .B0(n4093), .B1(n3843), .C0(n4252), 
        .C1(n3939), .Y(n1929) );
  OAI222XL U2840 ( .A0(n907), .A1(n3179), .B0(n4096), .B1(n3843), .C0(n4251), 
        .C1(n3940), .Y(n1928) );
  OAI222XL U2841 ( .A0(n908), .A1(n3179), .B0(n4099), .B1(n3842), .C0(n4250), 
        .C1(n3939), .Y(n1927) );
  OAI222XL U2842 ( .A0(n909), .A1(n3179), .B0(n4102), .B1(n3842), .C0(n4249), 
        .C1(n3940), .Y(n1926) );
  OAI222XL U2843 ( .A0(n910), .A1(n3179), .B0(n4105), .B1(n3842), .C0(n4248), 
        .C1(n3940), .Y(n1925) );
  OAI222XL U2844 ( .A0(n911), .A1(n3179), .B0(n4108), .B1(n3842), .C0(n4247), 
        .C1(n3940), .Y(n1924) );
  OAI222XL U2845 ( .A0(n912), .A1(n3179), .B0(n4111), .B1(n3842), .C0(n4246), 
        .C1(n3940), .Y(n1923) );
  OAI222XL U2846 ( .A0(n913), .A1(n3179), .B0(n4029), .B1(n3842), .C0(n4245), 
        .C1(n3940), .Y(n1922) );
  OAI222XL U2847 ( .A0(n914), .A1(n3179), .B0(n4031), .B1(n3842), .C0(n4244), 
        .C1(n3940), .Y(n1921) );
  OAI222XL U2848 ( .A0(n915), .A1(n3179), .B0(n4033), .B1(n3842), .C0(n4243), 
        .C1(n3940), .Y(n1920) );
  OAI222XL U2849 ( .A0(n916), .A1(n3179), .B0(n4035), .B1(n3842), .C0(n4242), 
        .C1(n3940), .Y(n1919) );
  OAI222XL U2850 ( .A0(n917), .A1(n3179), .B0(n4037), .B1(n3842), .C0(n4241), 
        .C1(n3940), .Y(n1918) );
  OAI222XL U2851 ( .A0(n918), .A1(n3179), .B0(n4039), .B1(n3842), .C0(n4240), 
        .C1(n3940), .Y(n1917) );
  OAI222XL U2852 ( .A0(n919), .A1(n3179), .B0(n4041), .B1(n3842), .C0(n4239), 
        .C1(n3940), .Y(n1916) );
  OAI222XL U2853 ( .A0(n1016), .A1(n3177), .B0(n4044), .B1(n3851), .C0(n4270), 
        .C1(n3951), .Y(n1819) );
  OAI222XL U2854 ( .A0(n1017), .A1(n3177), .B0(n4047), .B1(n3850), .C0(n4269), 
        .C1(n3952), .Y(n1818) );
  OAI222XL U2855 ( .A0(n1018), .A1(n3177), .B0(n4049), .B1(n327), .C0(n4268), 
        .C1(n3954), .Y(n1817) );
  OAI222XL U2856 ( .A0(n1019), .A1(n3177), .B0(n4051), .B1(n327), .C0(n4267), 
        .C1(n3953), .Y(n1816) );
  OAI222XL U2857 ( .A0(n1020), .A1(n3177), .B0(n4053), .B1(n327), .C0(n4266), 
        .C1(n3953), .Y(n1815) );
  OAI222XL U2858 ( .A0(n1021), .A1(n3177), .B0(n4055), .B1(n327), .C0(n4265), 
        .C1(n3952), .Y(n1814) );
  OAI222XL U2859 ( .A0(n1022), .A1(n3177), .B0(n4057), .B1(n327), .C0(n4264), 
        .C1(n3952), .Y(n1813) );
  OAI222XL U2860 ( .A0(n1023), .A1(n3177), .B0(n4059), .B1(n327), .C0(n4263), 
        .C1(n3952), .Y(n1812) );
  OAI222XL U2861 ( .A0(n1024), .A1(n3177), .B0(n4062), .B1(n3851), .C0(n4262), 
        .C1(n3952), .Y(n1811) );
  OAI222XL U2862 ( .A0(n1025), .A1(n3177), .B0(n4065), .B1(n3851), .C0(n4261), 
        .C1(n3952), .Y(n1810) );
  OAI222XL U2863 ( .A0(n1026), .A1(n3177), .B0(n4068), .B1(n3851), .C0(n4260), 
        .C1(n3952), .Y(n1809) );
  OAI222XL U2864 ( .A0(n1027), .A1(n3177), .B0(n4071), .B1(n3851), .C0(n4259), 
        .C1(n3952), .Y(n1808) );
  OAI222XL U2865 ( .A0(n1028), .A1(n3177), .B0(n4074), .B1(n3851), .C0(n4258), 
        .C1(n3952), .Y(n1807) );
  OAI222XL U2866 ( .A0(n1029), .A1(n3177), .B0(n4077), .B1(n3851), .C0(n4257), 
        .C1(n3952), .Y(n1806) );
  OAI222XL U2867 ( .A0(n1030), .A1(n3177), .B0(n4080), .B1(n3851), .C0(n4256), 
        .C1(n3952), .Y(n1805) );
  OAI222XL U2868 ( .A0(n1031), .A1(n3177), .B0(n4083), .B1(n3851), .C0(n4255), 
        .C1(n3952), .Y(n1804) );
  OAI222XL U2869 ( .A0(n1032), .A1(n3177), .B0(n4086), .B1(n3851), .C0(n4254), 
        .C1(n3952), .Y(n1803) );
  OAI222XL U2870 ( .A0(n1033), .A1(n3177), .B0(n4089), .B1(n3851), .C0(n4253), 
        .C1(n3952), .Y(n1802) );
  OAI222XL U2871 ( .A0(n1034), .A1(n3177), .B0(n4092), .B1(n3851), .C0(n4252), 
        .C1(n3952), .Y(n1801) );
  OAI222XL U2872 ( .A0(n1035), .A1(n3177), .B0(n4095), .B1(n3851), .C0(n4251), 
        .C1(n3953), .Y(n1800) );
  OAI222XL U2873 ( .A0(n1036), .A1(n3177), .B0(n4098), .B1(n3850), .C0(n4250), 
        .C1(n3952), .Y(n1799) );
  OAI222XL U2874 ( .A0(n1037), .A1(n3177), .B0(n4101), .B1(n3850), .C0(n4249), 
        .C1(n3953), .Y(n1798) );
  OAI222XL U2875 ( .A0(n1038), .A1(n3177), .B0(n4104), .B1(n3850), .C0(n4248), 
        .C1(n3953), .Y(n1797) );
  OAI222XL U2876 ( .A0(n1039), .A1(n3177), .B0(n4107), .B1(n3850), .C0(n4247), 
        .C1(n3953), .Y(n1796) );
  OAI222XL U2877 ( .A0(n1040), .A1(n3177), .B0(n4111), .B1(n3850), .C0(n4246), 
        .C1(n3953), .Y(n1795) );
  OAI222XL U2878 ( .A0(n1041), .A1(n3177), .B0(n4029), .B1(n3850), .C0(n4245), 
        .C1(n3953), .Y(n1794) );
  OAI222XL U2879 ( .A0(n1042), .A1(n3177), .B0(n4031), .B1(n3850), .C0(n4244), 
        .C1(n3953), .Y(n1793) );
  OAI222XL U2880 ( .A0(n1043), .A1(n3177), .B0(n4033), .B1(n3850), .C0(n4243), 
        .C1(n3953), .Y(n1792) );
  OAI222XL U2881 ( .A0(n1044), .A1(n3177), .B0(n4035), .B1(n3850), .C0(n4242), 
        .C1(n3953), .Y(n1791) );
  OAI222XL U2882 ( .A0(n1045), .A1(n3177), .B0(n4037), .B1(n3850), .C0(n4241), 
        .C1(n3953), .Y(n1790) );
  OAI222XL U2883 ( .A0(n1046), .A1(n3177), .B0(n4039), .B1(n3850), .C0(n4240), 
        .C1(n3953), .Y(n1789) );
  OAI222XL U2884 ( .A0(n1047), .A1(n3177), .B0(n4041), .B1(n3850), .C0(n4239), 
        .C1(n3953), .Y(n1788) );
  OAI222XL U2885 ( .A0(n1415), .A1(n4014), .B0(n4044), .B1(n4011), .C0(n4270), 
        .C1(n3860), .Y(n2715) );
  OAI222XL U2886 ( .A0(n1416), .A1(n4014), .B0(n4047), .B1(n4011), .C0(n4269), 
        .C1(n3864), .Y(n2714) );
  OAI222XL U2887 ( .A0(n1417), .A1(n4014), .B0(n4049), .B1(n4011), .C0(n4268), 
        .C1(n3861), .Y(n2713) );
  OAI222XL U2888 ( .A0(n1418), .A1(n4014), .B0(n4051), .B1(n4011), .C0(n4267), 
        .C1(n3865), .Y(n2712) );
  OAI222XL U2889 ( .A0(n1419), .A1(n4014), .B0(n4053), .B1(n4011), .C0(n4266), 
        .C1(n3858), .Y(n2711) );
  OAI222XL U2890 ( .A0(n1420), .A1(n4014), .B0(n4055), .B1(n4011), .C0(n4265), 
        .C1(n3865), .Y(n2710) );
  OAI222XL U2891 ( .A0(n1421), .A1(n4014), .B0(n4057), .B1(n4011), .C0(n4264), 
        .C1(n3861), .Y(n2709) );
  OAI222XL U2892 ( .A0(n1422), .A1(n4014), .B0(n4059), .B1(n4011), .C0(n4263), 
        .C1(n3858), .Y(n2708) );
  OAI222XL U2893 ( .A0(n1423), .A1(n4014), .B0(n4062), .B1(n4013), .C0(n4262), 
        .C1(n3865), .Y(n2707) );
  OAI222XL U2894 ( .A0(n1424), .A1(n4014), .B0(n4065), .B1(n4013), .C0(n4261), 
        .C1(n3861), .Y(n2706) );
  OAI222XL U2895 ( .A0(n1425), .A1(n4014), .B0(n4068), .B1(n4013), .C0(n4260), 
        .C1(n3858), .Y(n2705) );
  OAI222XL U2896 ( .A0(n1426), .A1(n4014), .B0(n4071), .B1(n4013), .C0(n4259), 
        .C1(n3864), .Y(n2704) );
  OAI222XL U2897 ( .A0(n1427), .A1(n4014), .B0(n4074), .B1(n4013), .C0(n4258), 
        .C1(n3862), .Y(n2703) );
  OAI222XL U2898 ( .A0(n1428), .A1(n4014), .B0(n4077), .B1(n4013), .C0(n4257), 
        .C1(n3863), .Y(n2702) );
  OAI222XL U2899 ( .A0(n1429), .A1(n4014), .B0(n4080), .B1(n4013), .C0(n4256), 
        .C1(n3862), .Y(n2701) );
  OAI222XL U2900 ( .A0(n1430), .A1(n4014), .B0(n4083), .B1(n4013), .C0(n4255), 
        .C1(n3863), .Y(n2700) );
  OAI222XL U2901 ( .A0(n1431), .A1(n4014), .B0(n4086), .B1(n4013), .C0(n4254), 
        .C1(n3862), .Y(n2699) );
  OAI222XL U2902 ( .A0(n1432), .A1(n4014), .B0(n4089), .B1(n4013), .C0(n4253), 
        .C1(n3863), .Y(n2698) );
  OAI222XL U2903 ( .A0(n1433), .A1(n4014), .B0(n4092), .B1(n4013), .C0(n4252), 
        .C1(n3862), .Y(n2697) );
  OAI222XL U2904 ( .A0(n1434), .A1(n4014), .B0(n4095), .B1(n4013), .C0(n4251), 
        .C1(n3862), .Y(n2696) );
  OAI222XL U2905 ( .A0(n1435), .A1(n4014), .B0(n4098), .B1(n4012), .C0(n4250), 
        .C1(n3862), .Y(n2695) );
  OAI222XL U2906 ( .A0(n1436), .A1(n4014), .B0(n4101), .B1(n4012), .C0(n4249), 
        .C1(n3862), .Y(n2694) );
  OAI222XL U2907 ( .A0(n1437), .A1(n4014), .B0(n4104), .B1(n4012), .C0(n4248), 
        .C1(n3862), .Y(n2693) );
  OAI222XL U2908 ( .A0(n1438), .A1(n4014), .B0(n4107), .B1(n4012), .C0(n4247), 
        .C1(n3862), .Y(n2692) );
  OAI222XL U2909 ( .A0(n1439), .A1(n4014), .B0(n4110), .B1(n4012), .C0(n4246), 
        .C1(n3862), .Y(n2691) );
  OAI222XL U2910 ( .A0(n1440), .A1(n4014), .B0(n4028), .B1(n4012), .C0(n4245), 
        .C1(n3862), .Y(n2690) );
  OAI222XL U2911 ( .A0(n1441), .A1(n4014), .B0(n4030), .B1(n4012), .C0(n4244), 
        .C1(n3862), .Y(n2689) );
  OAI222XL U2912 ( .A0(n1442), .A1(n4014), .B0(n4032), .B1(n4012), .C0(n4243), 
        .C1(n3862), .Y(n2688) );
  OAI222XL U2913 ( .A0(n1443), .A1(n4014), .B0(n4034), .B1(n4012), .C0(n4242), 
        .C1(n3862), .Y(n2687) );
  OAI222XL U2914 ( .A0(n1444), .A1(n4014), .B0(n4036), .B1(n4012), .C0(n4241), 
        .C1(n3862), .Y(n2686) );
  OAI222XL U2915 ( .A0(n1445), .A1(n4014), .B0(n4038), .B1(n4012), .C0(n4240), 
        .C1(n3862), .Y(n2685) );
  OAI222XL U2916 ( .A0(n1446), .A1(n4014), .B0(n4040), .B1(n4012), .C0(n4239), 
        .C1(n3862), .Y(n2684) );
  OAI222XL U2917 ( .A0(n1543), .A1(n4025), .B0(n4044), .B1(n4022), .C0(n4270), 
        .C1(n3874), .Y(n2587) );
  OAI222XL U2918 ( .A0(n1544), .A1(n4025), .B0(n4047), .B1(n4022), .C0(n4269), 
        .C1(n3874), .Y(n2586) );
  OAI222XL U2919 ( .A0(n1545), .A1(n4025), .B0(n4049), .B1(n4022), .C0(n4268), 
        .C1(n3874), .Y(n2585) );
  OAI222XL U2920 ( .A0(n1546), .A1(n4025), .B0(n4051), .B1(n4022), .C0(n4267), 
        .C1(n3874), .Y(n2584) );
  OAI222XL U2921 ( .A0(n1547), .A1(n4025), .B0(n4053), .B1(n4022), .C0(n4266), 
        .C1(n3875), .Y(n2583) );
  OAI222XL U2922 ( .A0(n1548), .A1(n4025), .B0(n4055), .B1(n4022), .C0(n4265), 
        .C1(n3875), .Y(n2582) );
  OAI222XL U2923 ( .A0(n1549), .A1(n4025), .B0(n4057), .B1(n4022), .C0(n4264), 
        .C1(n3875), .Y(n2581) );
  OAI222XL U2924 ( .A0(n1550), .A1(n4025), .B0(n4059), .B1(n4022), .C0(n4263), 
        .C1(n3875), .Y(n2580) );
  OAI222XL U2925 ( .A0(n1551), .A1(n4025), .B0(n4062), .B1(n4024), .C0(n4262), 
        .C1(n3875), .Y(n2579) );
  OAI222XL U2926 ( .A0(n1552), .A1(n4025), .B0(n4065), .B1(n4024), .C0(n4261), 
        .C1(n3875), .Y(n2578) );
  OAI222XL U2927 ( .A0(n1553), .A1(n4025), .B0(n4068), .B1(n4024), .C0(n4260), 
        .C1(n3875), .Y(n2577) );
  OAI222XL U2928 ( .A0(n1554), .A1(n4025), .B0(n4071), .B1(n4024), .C0(n4259), 
        .C1(n3875), .Y(n2576) );
  OAI222XL U2929 ( .A0(n1555), .A1(n4025), .B0(n4074), .B1(n4024), .C0(n4258), 
        .C1(n3875), .Y(n2575) );
  OAI222XL U2930 ( .A0(n1556), .A1(n4025), .B0(n4077), .B1(n4024), .C0(n4257), 
        .C1(n3875), .Y(n2574) );
  OAI222XL U2931 ( .A0(n1557), .A1(n4025), .B0(n4080), .B1(n4024), .C0(n4256), 
        .C1(n3875), .Y(n2573) );
  OAI222XL U2932 ( .A0(n1558), .A1(n4025), .B0(n4083), .B1(n4024), .C0(n4255), 
        .C1(n3875), .Y(n2572) );
  OAI222XL U2933 ( .A0(n1559), .A1(n4025), .B0(n4086), .B1(n4024), .C0(n4254), 
        .C1(n3875), .Y(n2571) );
  OAI222XL U2934 ( .A0(n1560), .A1(n4025), .B0(n4089), .B1(n4024), .C0(n4253), 
        .C1(n3875), .Y(n2570) );
  OAI222XL U2935 ( .A0(n1561), .A1(n4025), .B0(n4092), .B1(n4024), .C0(n4252), 
        .C1(n3875), .Y(n2569) );
  OAI222XL U2936 ( .A0(n1562), .A1(n4025), .B0(n4095), .B1(n4024), .C0(n4251), 
        .C1(n3875), .Y(n2568) );
  OAI222XL U2937 ( .A0(n1563), .A1(n4025), .B0(n4098), .B1(n4023), .C0(n4250), 
        .C1(n3876), .Y(n2567) );
  OAI222XL U2938 ( .A0(n1564), .A1(n4025), .B0(n4101), .B1(n4023), .C0(n4249), 
        .C1(n3876), .Y(n2566) );
  OAI222XL U2939 ( .A0(n1565), .A1(n4025), .B0(n4104), .B1(n4023), .C0(n4248), 
        .C1(n3876), .Y(n2565) );
  OAI222XL U2940 ( .A0(n1566), .A1(n4025), .B0(n4107), .B1(n4023), .C0(n4247), 
        .C1(n3876), .Y(n2564) );
  OAI222XL U2941 ( .A0(n1567), .A1(n4025), .B0(n4110), .B1(n4023), .C0(n4246), 
        .C1(n3876), .Y(n2563) );
  OAI222XL U2942 ( .A0(n1568), .A1(n4025), .B0(n4029), .B1(n4023), .C0(n3876), 
        .C1(n4245), .Y(n2562) );
  OAI222XL U2943 ( .A0(n1569), .A1(n4025), .B0(n4031), .B1(n4023), .C0(n3876), 
        .C1(n4244), .Y(n2561) );
  OAI222XL U2944 ( .A0(n1570), .A1(n4025), .B0(n4033), .B1(n4023), .C0(n3876), 
        .C1(n4243), .Y(n2560) );
  OAI222XL U2945 ( .A0(n1571), .A1(n4025), .B0(n4035), .B1(n4023), .C0(n3876), 
        .C1(n4242), .Y(n2559) );
  OAI222XL U2946 ( .A0(n1572), .A1(n4025), .B0(n4037), .B1(n4023), .C0(n3876), 
        .C1(n4241), .Y(n2558) );
  OAI222XL U2947 ( .A0(n1573), .A1(n4025), .B0(n4039), .B1(n4023), .C0(n3876), 
        .C1(n4240), .Y(n2557) );
  OAI222XL U2948 ( .A0(n1574), .A1(n4025), .B0(n4041), .B1(n4023), .C0(n3876), 
        .C1(n4239), .Y(n2556) );
  OAI222XL U2949 ( .A0(n408), .A1(n3202), .B0(n4043), .B1(n3813), .C0(n3886), 
        .C1(n4238), .Y(n2427) );
  OAI222XL U2950 ( .A0(n409), .A1(n3202), .B0(n4046), .B1(n3812), .C0(n3887), 
        .C1(n4237), .Y(n2426) );
  OAI222XL U2951 ( .A0(n410), .A1(n3202), .B0(n4050), .B1(n367), .C0(n3885), 
        .C1(n4236), .Y(n2425) );
  OAI222XL U2952 ( .A0(n411), .A1(n3202), .B0(n4052), .B1(n367), .C0(n3885), 
        .C1(n4235), .Y(n2424) );
  OAI222XL U2953 ( .A0(n412), .A1(n3202), .B0(n4054), .B1(n367), .C0(n3885), 
        .C1(n4234), .Y(n2423) );
  OAI222XL U2954 ( .A0(n413), .A1(n3202), .B0(n4056), .B1(n367), .C0(n3885), 
        .C1(n4233), .Y(n2422) );
  OAI222XL U2955 ( .A0(n414), .A1(n3202), .B0(n4058), .B1(n367), .C0(n3890), 
        .C1(n4232), .Y(n2421) );
  OAI222XL U2956 ( .A0(n415), .A1(n3202), .B0(n4060), .B1(n367), .C0(n3886), 
        .C1(n4231), .Y(n2420) );
  OAI222XL U2957 ( .A0(n416), .A1(n3202), .B0(n4061), .B1(n3813), .C0(n3885), 
        .C1(n4230), .Y(n2419) );
  OAI222XL U2958 ( .A0(n417), .A1(n3202), .B0(n4064), .B1(n3813), .C0(n3888), 
        .C1(n4229), .Y(n2418) );
  OAI222XL U2959 ( .A0(n418), .A1(n3202), .B0(n4067), .B1(n3813), .C0(n3885), 
        .C1(n4228), .Y(n2417) );
  OAI222XL U2960 ( .A0(n419), .A1(n3202), .B0(n4070), .B1(n3813), .C0(n3886), 
        .C1(n4227), .Y(n2416) );
  OAI222XL U2961 ( .A0(n420), .A1(n3202), .B0(n4073), .B1(n3813), .C0(n3890), 
        .C1(n4226), .Y(n2415) );
  OAI222XL U2962 ( .A0(n421), .A1(n3202), .B0(n4076), .B1(n3813), .C0(n3886), 
        .C1(n4225), .Y(n2414) );
  OAI222XL U2963 ( .A0(n422), .A1(n3202), .B0(n4079), .B1(n3813), .C0(n3886), 
        .C1(n4224), .Y(n2413) );
  OAI222XL U2964 ( .A0(n423), .A1(n3202), .B0(n4082), .B1(n3813), .C0(n3887), 
        .C1(n4223), .Y(n2412) );
  OAI222XL U2965 ( .A0(n424), .A1(n3202), .B0(n4085), .B1(n3813), .C0(n3888), 
        .C1(n4222), .Y(n2411) );
  OAI222XL U2966 ( .A0(n425), .A1(n3202), .B0(n4088), .B1(n3813), .C0(n3886), 
        .C1(n4221), .Y(n2410) );
  OAI222XL U2967 ( .A0(n426), .A1(n3202), .B0(n4091), .B1(n3813), .C0(n3890), 
        .C1(n4220), .Y(n2409) );
  OAI222XL U2968 ( .A0(n427), .A1(n3202), .B0(n4094), .B1(n3813), .C0(n3886), 
        .C1(n4219), .Y(n2408) );
  OAI222XL U2969 ( .A0(n428), .A1(n3202), .B0(n4097), .B1(n3812), .C0(n3886), 
        .C1(n4218), .Y(n2407) );
  OAI222XL U2970 ( .A0(n429), .A1(n3202), .B0(n4100), .B1(n3812), .C0(n3886), 
        .C1(n4217), .Y(n2406) );
  OAI222XL U2971 ( .A0(n430), .A1(n3202), .B0(n4103), .B1(n3812), .C0(n3887), 
        .C1(n4216), .Y(n2405) );
  OAI222XL U2972 ( .A0(n431), .A1(n3202), .B0(n4106), .B1(n3812), .C0(n3886), 
        .C1(n4215), .Y(n2404) );
  OAI222XL U2973 ( .A0(n432), .A1(n3202), .B0(n4111), .B1(n3812), .C0(n3888), 
        .C1(n4214), .Y(n2403) );
  OAI222XL U2974 ( .A0(n433), .A1(n3202), .B0(n4028), .B1(n3812), .C0(n3885), 
        .C1(n4213), .Y(n2402) );
  OAI222XL U2975 ( .A0(n434), .A1(n3202), .B0(n4030), .B1(n3812), .C0(n3886), 
        .C1(n4212), .Y(n2401) );
  OAI222XL U2976 ( .A0(n435), .A1(n3202), .B0(n4032), .B1(n3812), .C0(n3886), 
        .C1(n4211), .Y(n2400) );
  OAI222XL U2977 ( .A0(n436), .A1(n3202), .B0(n4034), .B1(n3812), .C0(n3885), 
        .C1(n4210), .Y(n2399) );
  OAI222XL U2978 ( .A0(n437), .A1(n3202), .B0(n4036), .B1(n3812), .C0(n3887), 
        .C1(n4209), .Y(n2398) );
  OAI222XL U2979 ( .A0(n438), .A1(n3202), .B0(n4038), .B1(n3812), .C0(n3885), 
        .C1(n4208), .Y(n2397) );
  OAI222XL U2980 ( .A0(n439), .A1(n3202), .B0(n4040), .B1(n3812), .C0(n3885), 
        .C1(n4207), .Y(n2396) );
  OAI222XL U2981 ( .A0(n536), .A1(n3192), .B0(n4043), .B1(n3821), .C0(n4238), 
        .C1(n3901), .Y(n2299) );
  OAI222XL U2982 ( .A0(n537), .A1(n3192), .B0(n4046), .B1(n3820), .C0(n4237), 
        .C1(n3901), .Y(n2298) );
  OAI222XL U2983 ( .A0(n538), .A1(n3192), .B0(n4049), .B1(n357), .C0(n4236), 
        .C1(n3901), .Y(n2297) );
  OAI222XL U2984 ( .A0(n539), .A1(n3192), .B0(n4051), .B1(n357), .C0(n4235), 
        .C1(n3902), .Y(n2296) );
  OAI222XL U2985 ( .A0(n540), .A1(n3192), .B0(n4053), .B1(n357), .C0(n4234), 
        .C1(n3902), .Y(n2295) );
  OAI222XL U2986 ( .A0(n541), .A1(n3192), .B0(n4055), .B1(n357), .C0(n4233), 
        .C1(n3902), .Y(n2294) );
  OAI222XL U2987 ( .A0(n542), .A1(n3192), .B0(n4057), .B1(n357), .C0(n4232), 
        .C1(n3902), .Y(n2293) );
  OAI222XL U2988 ( .A0(n543), .A1(n3192), .B0(n4059), .B1(n357), .C0(n4231), 
        .C1(n3902), .Y(n2292) );
  OAI222XL U2989 ( .A0(n544), .A1(n3192), .B0(n4061), .B1(n3821), .C0(n4230), 
        .C1(n3902), .Y(n2291) );
  OAI222XL U2990 ( .A0(n545), .A1(n3192), .B0(n4064), .B1(n3821), .C0(n4229), 
        .C1(n3902), .Y(n2290) );
  OAI222XL U2991 ( .A0(n546), .A1(n3192), .B0(n4067), .B1(n3821), .C0(n4228), 
        .C1(n3902), .Y(n2289) );
  OAI222XL U2992 ( .A0(n547), .A1(n3192), .B0(n4070), .B1(n3821), .C0(n4227), 
        .C1(n3902), .Y(n2288) );
  OAI222XL U2993 ( .A0(n548), .A1(n3192), .B0(n4073), .B1(n3821), .C0(n4226), 
        .C1(n3902), .Y(n2287) );
  OAI222XL U2994 ( .A0(n549), .A1(n3192), .B0(n4076), .B1(n3821), .C0(n4225), 
        .C1(n3902), .Y(n2286) );
  OAI222XL U2995 ( .A0(n550), .A1(n3192), .B0(n4079), .B1(n3821), .C0(n4224), 
        .C1(n3902), .Y(n2285) );
  OAI222XL U2996 ( .A0(n551), .A1(n3192), .B0(n4082), .B1(n3821), .C0(n4223), 
        .C1(n3902), .Y(n2284) );
  OAI222XL U2997 ( .A0(n552), .A1(n3192), .B0(n4085), .B1(n3821), .C0(n4222), 
        .C1(n3902), .Y(n2283) );
  OAI222XL U2998 ( .A0(n553), .A1(n3192), .B0(n4088), .B1(n3821), .C0(n4221), 
        .C1(n3902), .Y(n2282) );
  OAI222XL U2999 ( .A0(n554), .A1(n3192), .B0(n4091), .B1(n3821), .C0(n4220), 
        .C1(n3902), .Y(n2281) );
  OAI222XL U3000 ( .A0(n555), .A1(n3192), .B0(n4094), .B1(n3821), .C0(n4219), 
        .C1(n3903), .Y(n2280) );
  OAI222XL U3001 ( .A0(n556), .A1(n3192), .B0(n4097), .B1(n3820), .C0(n4218), 
        .C1(n3903), .Y(n2279) );
  OAI222XL U3002 ( .A0(n557), .A1(n3192), .B0(n4100), .B1(n3820), .C0(n4217), 
        .C1(n3903), .Y(n2278) );
  OAI222XL U3003 ( .A0(n558), .A1(n3192), .B0(n4103), .B1(n3820), .C0(n4216), 
        .C1(n3903), .Y(n2277) );
  OAI222XL U3004 ( .A0(n559), .A1(n3192), .B0(n4106), .B1(n3820), .C0(n4215), 
        .C1(n3903), .Y(n2276) );
  OAI222XL U3005 ( .A0(n560), .A1(n3192), .B0(n4110), .B1(n3820), .C0(n4214), 
        .C1(n3903), .Y(n2275) );
  OAI222XL U3006 ( .A0(n561), .A1(n3192), .B0(n4028), .B1(n3820), .C0(n4213), 
        .C1(n3903), .Y(n2274) );
  OAI222XL U3007 ( .A0(n562), .A1(n3192), .B0(n4030), .B1(n3820), .C0(n4212), 
        .C1(n3903), .Y(n2273) );
  OAI222XL U3008 ( .A0(n563), .A1(n3192), .B0(n4032), .B1(n3820), .C0(n4211), 
        .C1(n3903), .Y(n2272) );
  OAI222XL U3009 ( .A0(n564), .A1(n3192), .B0(n4034), .B1(n3820), .C0(n4210), 
        .C1(n3903), .Y(n2271) );
  OAI222XL U3010 ( .A0(n565), .A1(n3192), .B0(n4036), .B1(n3820), .C0(n4209), 
        .C1(n3903), .Y(n2270) );
  OAI222XL U3011 ( .A0(n566), .A1(n3192), .B0(n4038), .B1(n3820), .C0(n4208), 
        .C1(n3903), .Y(n2269) );
  OAI222XL U3012 ( .A0(n567), .A1(n3192), .B0(n4040), .B1(n3820), .C0(n4207), 
        .C1(n3903), .Y(n2268) );
  OAI222XL U3013 ( .A0(n664), .A1(n3191), .B0(n4045), .B1(n3829), .C0(n4238), 
        .C1(n3914), .Y(n2171) );
  OAI222XL U3014 ( .A0(n665), .A1(n3191), .B0(n4048), .B1(n3828), .C0(n4237), 
        .C1(n3914), .Y(n2170) );
  OAI222XL U3015 ( .A0(n666), .A1(n3191), .B0(n4050), .B1(n349), .C0(n4236), 
        .C1(n3914), .Y(n2169) );
  OAI222XL U3016 ( .A0(n667), .A1(n3191), .B0(n4052), .B1(n349), .C0(n4235), 
        .C1(n3915), .Y(n2168) );
  OAI222XL U3017 ( .A0(n668), .A1(n3191), .B0(n4054), .B1(n349), .C0(n4234), 
        .C1(n3915), .Y(n2167) );
  OAI222XL U3018 ( .A0(n669), .A1(n3191), .B0(n4056), .B1(n349), .C0(n4233), 
        .C1(n3915), .Y(n2166) );
  OAI222XL U3019 ( .A0(n670), .A1(n3191), .B0(n4058), .B1(n349), .C0(n4232), 
        .C1(n3915), .Y(n2165) );
  OAI222XL U3020 ( .A0(n671), .A1(n3191), .B0(n4060), .B1(n349), .C0(n4231), 
        .C1(n3915), .Y(n2164) );
  OAI222XL U3021 ( .A0(n672), .A1(n3191), .B0(n4063), .B1(n3829), .C0(n4230), 
        .C1(n3915), .Y(n2163) );
  OAI222XL U3022 ( .A0(n673), .A1(n3191), .B0(n4066), .B1(n3829), .C0(n4229), 
        .C1(n3915), .Y(n2162) );
  OAI222XL U3023 ( .A0(n674), .A1(n3191), .B0(n4069), .B1(n3829), .C0(n4228), 
        .C1(n3915), .Y(n2161) );
  OAI222XL U3024 ( .A0(n675), .A1(n3191), .B0(n4072), .B1(n3829), .C0(n4227), 
        .C1(n3915), .Y(n2160) );
  OAI222XL U3025 ( .A0(n676), .A1(n3191), .B0(n4075), .B1(n3829), .C0(n4226), 
        .C1(n3915), .Y(n2159) );
  OAI222XL U3026 ( .A0(n677), .A1(n3191), .B0(n4078), .B1(n3829), .C0(n4225), 
        .C1(n3915), .Y(n2158) );
  OAI222XL U3027 ( .A0(n678), .A1(n3191), .B0(n4081), .B1(n3829), .C0(n4224), 
        .C1(n3915), .Y(n2157) );
  OAI222XL U3028 ( .A0(n679), .A1(n3191), .B0(n4084), .B1(n3829), .C0(n4223), 
        .C1(n3915), .Y(n2156) );
  OAI222XL U3029 ( .A0(n680), .A1(n3191), .B0(n4087), .B1(n3829), .C0(n4222), 
        .C1(n3915), .Y(n2155) );
  OAI222XL U3030 ( .A0(n681), .A1(n3191), .B0(n4090), .B1(n3829), .C0(n4221), 
        .C1(n3915), .Y(n2154) );
  OAI222XL U3031 ( .A0(n682), .A1(n3191), .B0(n4093), .B1(n3829), .C0(n4220), 
        .C1(n3915), .Y(n2153) );
  OAI222XL U3032 ( .A0(n683), .A1(n3191), .B0(n4096), .B1(n3829), .C0(n4219), 
        .C1(n3916), .Y(n2152) );
  OAI222XL U3033 ( .A0(n684), .A1(n3191), .B0(n4099), .B1(n3828), .C0(n4218), 
        .C1(n3916), .Y(n2151) );
  OAI222XL U3034 ( .A0(n685), .A1(n3191), .B0(n4102), .B1(n3828), .C0(n4217), 
        .C1(n3916), .Y(n2150) );
  OAI222XL U3035 ( .A0(n686), .A1(n3191), .B0(n4105), .B1(n3828), .C0(n4216), 
        .C1(n3916), .Y(n2149) );
  OAI222XL U3036 ( .A0(n687), .A1(n3191), .B0(n4108), .B1(n3828), .C0(n4215), 
        .C1(n3916), .Y(n2148) );
  OAI222XL U3037 ( .A0(n688), .A1(n3191), .B0(n4111), .B1(n3828), .C0(n4214), 
        .C1(n3916), .Y(n2147) );
  OAI222XL U3038 ( .A0(n689), .A1(n3191), .B0(n4028), .B1(n3828), .C0(n4213), 
        .C1(n3916), .Y(n2146) );
  OAI222XL U3039 ( .A0(n690), .A1(n3191), .B0(n4030), .B1(n3828), .C0(n4212), 
        .C1(n3916), .Y(n2145) );
  OAI222XL U3040 ( .A0(n691), .A1(n3191), .B0(n4032), .B1(n3828), .C0(n4211), 
        .C1(n3916), .Y(n2144) );
  OAI222XL U3041 ( .A0(n692), .A1(n3191), .B0(n4034), .B1(n3828), .C0(n4210), 
        .C1(n3916), .Y(n2143) );
  OAI222XL U3042 ( .A0(n693), .A1(n3191), .B0(n4036), .B1(n3828), .C0(n4209), 
        .C1(n3916), .Y(n2142) );
  OAI222XL U3043 ( .A0(n694), .A1(n3191), .B0(n4038), .B1(n3828), .C0(n4208), 
        .C1(n3916), .Y(n2141) );
  OAI222XL U3044 ( .A0(n695), .A1(n3191), .B0(n4040), .B1(n3828), .C0(n4207), 
        .C1(n3916), .Y(n2140) );
  OAI222XL U3045 ( .A0(n792), .A1(n3195), .B0(n4045), .B1(n3837), .C0(n4238), 
        .C1(n3927), .Y(n2043) );
  OAI222XL U3046 ( .A0(n793), .A1(n3195), .B0(n4048), .B1(n3836), .C0(n4237), 
        .C1(n3927), .Y(n2042) );
  OAI222XL U3047 ( .A0(n794), .A1(n3195), .B0(n4050), .B1(n341), .C0(n4236), 
        .C1(n3927), .Y(n2041) );
  OAI222XL U3048 ( .A0(n795), .A1(n3195), .B0(n4052), .B1(n341), .C0(n4235), 
        .C1(n3928), .Y(n2040) );
  OAI222XL U3049 ( .A0(n796), .A1(n3195), .B0(n4054), .B1(n341), .C0(n4234), 
        .C1(n3928), .Y(n2039) );
  OAI222XL U3050 ( .A0(n797), .A1(n3195), .B0(n4056), .B1(n341), .C0(n4233), 
        .C1(n3928), .Y(n2038) );
  OAI222XL U3051 ( .A0(n798), .A1(n3195), .B0(n4058), .B1(n341), .C0(n4232), 
        .C1(n3928), .Y(n2037) );
  OAI222XL U3052 ( .A0(n799), .A1(n3195), .B0(n4060), .B1(n341), .C0(n4231), 
        .C1(n3928), .Y(n2036) );
  OAI222XL U3053 ( .A0(n800), .A1(n3195), .B0(n4063), .B1(n3837), .C0(n4230), 
        .C1(n3928), .Y(n2035) );
  OAI222XL U3054 ( .A0(n801), .A1(n3195), .B0(n4066), .B1(n3837), .C0(n4229), 
        .C1(n3928), .Y(n2034) );
  OAI222XL U3055 ( .A0(n802), .A1(n3195), .B0(n4069), .B1(n3837), .C0(n4228), 
        .C1(n3928), .Y(n2033) );
  OAI222XL U3056 ( .A0(n803), .A1(n3195), .B0(n4072), .B1(n3837), .C0(n4227), 
        .C1(n3928), .Y(n2032) );
  OAI222XL U3057 ( .A0(n804), .A1(n3195), .B0(n4075), .B1(n3837), .C0(n4226), 
        .C1(n3928), .Y(n2031) );
  OAI222XL U3058 ( .A0(n805), .A1(n3195), .B0(n4078), .B1(n3837), .C0(n4225), 
        .C1(n3928), .Y(n2030) );
  OAI222XL U3059 ( .A0(n806), .A1(n3195), .B0(n4081), .B1(n3837), .C0(n4224), 
        .C1(n3928), .Y(n2029) );
  OAI222XL U3060 ( .A0(n807), .A1(n3195), .B0(n4084), .B1(n3837), .C0(n4223), 
        .C1(n3928), .Y(n2028) );
  OAI222XL U3061 ( .A0(n808), .A1(n3195), .B0(n4087), .B1(n3837), .C0(n4222), 
        .C1(n3928), .Y(n2027) );
  OAI222XL U3062 ( .A0(n809), .A1(n3195), .B0(n4090), .B1(n3837), .C0(n4221), 
        .C1(n3928), .Y(n2026) );
  OAI222XL U3063 ( .A0(n810), .A1(n3195), .B0(n4093), .B1(n3837), .C0(n4220), 
        .C1(n3928), .Y(n2025) );
  OAI222XL U3064 ( .A0(n811), .A1(n3195), .B0(n4096), .B1(n3837), .C0(n4219), 
        .C1(n3929), .Y(n2024) );
  OAI222XL U3065 ( .A0(n812), .A1(n3195), .B0(n4099), .B1(n3836), .C0(n4218), 
        .C1(n3929), .Y(n2023) );
  OAI222XL U3066 ( .A0(n813), .A1(n3195), .B0(n4102), .B1(n3836), .C0(n4217), 
        .C1(n3929), .Y(n2022) );
  OAI222XL U3067 ( .A0(n814), .A1(n3195), .B0(n4105), .B1(n3836), .C0(n4216), 
        .C1(n3929), .Y(n2021) );
  OAI222XL U3068 ( .A0(n815), .A1(n3195), .B0(n4108), .B1(n3836), .C0(n4215), 
        .C1(n3929), .Y(n2020) );
  OAI222XL U3069 ( .A0(n816), .A1(n3195), .B0(n4111), .B1(n3836), .C0(n4214), 
        .C1(n3929), .Y(n2019) );
  OAI222XL U3070 ( .A0(n817), .A1(n3195), .B0(n4029), .B1(n3836), .C0(n4213), 
        .C1(n3929), .Y(n2018) );
  OAI222XL U3071 ( .A0(n818), .A1(n3195), .B0(n4031), .B1(n3836), .C0(n4212), 
        .C1(n3929), .Y(n2017) );
  OAI222XL U3072 ( .A0(n819), .A1(n3195), .B0(n4033), .B1(n3836), .C0(n4211), 
        .C1(n3929), .Y(n2016) );
  OAI222XL U3073 ( .A0(n820), .A1(n3195), .B0(n4035), .B1(n3836), .C0(n4210), 
        .C1(n3929), .Y(n2015) );
  OAI222XL U3074 ( .A0(n821), .A1(n3195), .B0(n4037), .B1(n3836), .C0(n4209), 
        .C1(n3929), .Y(n2014) );
  OAI222XL U3075 ( .A0(n822), .A1(n3195), .B0(n4039), .B1(n3836), .C0(n4208), 
        .C1(n3929), .Y(n2013) );
  OAI222XL U3076 ( .A0(n823), .A1(n3195), .B0(n4041), .B1(n3836), .C0(n4207), 
        .C1(n3929), .Y(n2012) );
  OAI222XL U3077 ( .A0(n920), .A1(n3194), .B0(n4045), .B1(n3845), .C0(n4238), 
        .C1(n3940), .Y(n1915) );
  OAI222XL U3078 ( .A0(n921), .A1(n3194), .B0(n4048), .B1(n3844), .C0(n4237), 
        .C1(n3940), .Y(n1914) );
  OAI222XL U3079 ( .A0(n922), .A1(n3194), .B0(n4050), .B1(n333), .C0(n4236), 
        .C1(n3940), .Y(n1913) );
  OAI222XL U3080 ( .A0(n923), .A1(n3194), .B0(n4052), .B1(n333), .C0(n4235), 
        .C1(n3941), .Y(n1912) );
  OAI222XL U3081 ( .A0(n924), .A1(n3194), .B0(n4054), .B1(n333), .C0(n4234), 
        .C1(n3941), .Y(n1911) );
  OAI222XL U3082 ( .A0(n925), .A1(n3194), .B0(n4056), .B1(n333), .C0(n4233), 
        .C1(n3941), .Y(n1910) );
  OAI222XL U3083 ( .A0(n926), .A1(n3194), .B0(n4058), .B1(n333), .C0(n4232), 
        .C1(n3941), .Y(n1909) );
  OAI222XL U3084 ( .A0(n927), .A1(n3194), .B0(n4060), .B1(n333), .C0(n4231), 
        .C1(n3941), .Y(n1908) );
  OAI222XL U3085 ( .A0(n928), .A1(n3194), .B0(n4063), .B1(n3845), .C0(n4230), 
        .C1(n3941), .Y(n1907) );
  OAI222XL U3086 ( .A0(n929), .A1(n3194), .B0(n4066), .B1(n3845), .C0(n4229), 
        .C1(n3941), .Y(n1906) );
  OAI222XL U3087 ( .A0(n930), .A1(n3194), .B0(n4069), .B1(n3845), .C0(n4228), 
        .C1(n3941), .Y(n1905) );
  OAI222XL U3088 ( .A0(n931), .A1(n3194), .B0(n4072), .B1(n3845), .C0(n4227), 
        .C1(n3941), .Y(n1904) );
  OAI222XL U3089 ( .A0(n932), .A1(n3194), .B0(n4075), .B1(n3845), .C0(n4226), 
        .C1(n3941), .Y(n1903) );
  OAI222XL U3090 ( .A0(n933), .A1(n3194), .B0(n4078), .B1(n3845), .C0(n4225), 
        .C1(n3941), .Y(n1902) );
  OAI222XL U3091 ( .A0(n934), .A1(n3194), .B0(n4081), .B1(n3845), .C0(n4224), 
        .C1(n3941), .Y(n1901) );
  OAI222XL U3092 ( .A0(n935), .A1(n3194), .B0(n4084), .B1(n3845), .C0(n4223), 
        .C1(n3941), .Y(n1900) );
  OAI222XL U3093 ( .A0(n936), .A1(n3194), .B0(n4087), .B1(n3845), .C0(n4222), 
        .C1(n3941), .Y(n1899) );
  OAI222XL U3094 ( .A0(n937), .A1(n3194), .B0(n4090), .B1(n3845), .C0(n4221), 
        .C1(n3941), .Y(n1898) );
  OAI222XL U3095 ( .A0(n938), .A1(n3194), .B0(n4093), .B1(n3845), .C0(n4220), 
        .C1(n3941), .Y(n1897) );
  OAI222XL U3096 ( .A0(n939), .A1(n3194), .B0(n4096), .B1(n3845), .C0(n4219), 
        .C1(n3942), .Y(n1896) );
  OAI222XL U3097 ( .A0(n940), .A1(n3194), .B0(n4099), .B1(n3844), .C0(n4218), 
        .C1(n3942), .Y(n1895) );
  OAI222XL U3098 ( .A0(n941), .A1(n3194), .B0(n4102), .B1(n3844), .C0(n4217), 
        .C1(n3942), .Y(n1894) );
  OAI222XL U3099 ( .A0(n942), .A1(n3194), .B0(n4105), .B1(n3844), .C0(n4216), 
        .C1(n3942), .Y(n1893) );
  OAI222XL U3100 ( .A0(n943), .A1(n3194), .B0(n4108), .B1(n3844), .C0(n4215), 
        .C1(n3942), .Y(n1892) );
  OAI222XL U3101 ( .A0(n944), .A1(n3194), .B0(n4111), .B1(n3844), .C0(n4214), 
        .C1(n3942), .Y(n1891) );
  OAI222XL U3102 ( .A0(n945), .A1(n3194), .B0(n4029), .B1(n3844), .C0(n4213), 
        .C1(n3942), .Y(n1890) );
  OAI222XL U3103 ( .A0(n946), .A1(n3194), .B0(n4031), .B1(n3844), .C0(n4212), 
        .C1(n3942), .Y(n1889) );
  OAI222XL U3104 ( .A0(n947), .A1(n3194), .B0(n4033), .B1(n3844), .C0(n4211), 
        .C1(n3942), .Y(n1888) );
  OAI222XL U3105 ( .A0(n948), .A1(n3194), .B0(n4035), .B1(n3844), .C0(n4210), 
        .C1(n3942), .Y(n1887) );
  OAI222XL U3106 ( .A0(n949), .A1(n3194), .B0(n4037), .B1(n3844), .C0(n4209), 
        .C1(n3942), .Y(n1886) );
  OAI222XL U3107 ( .A0(n950), .A1(n3194), .B0(n4039), .B1(n3844), .C0(n4208), 
        .C1(n3942), .Y(n1885) );
  OAI222XL U3108 ( .A0(n951), .A1(n3194), .B0(n4041), .B1(n3844), .C0(n4207), 
        .C1(n3942), .Y(n1884) );
  OAI222XL U3109 ( .A0(n1048), .A1(n3193), .B0(n4044), .B1(n3853), .C0(n4238), 
        .C1(n3953), .Y(n1787) );
  OAI222XL U3110 ( .A0(n1049), .A1(n3193), .B0(n4047), .B1(n3852), .C0(n4237), 
        .C1(n3953), .Y(n1786) );
  OAI222XL U3111 ( .A0(n1050), .A1(n3193), .B0(n4049), .B1(n325), .C0(n4236), 
        .C1(n3953), .Y(n1785) );
  OAI222XL U3112 ( .A0(n1051), .A1(n3193), .B0(n4051), .B1(n325), .C0(n4235), 
        .C1(n3954), .Y(n1784) );
  OAI222XL U3113 ( .A0(n1052), .A1(n3193), .B0(n4053), .B1(n325), .C0(n4234), 
        .C1(n3954), .Y(n1783) );
  OAI222XL U3114 ( .A0(n1053), .A1(n3193), .B0(n4055), .B1(n325), .C0(n4233), 
        .C1(n3954), .Y(n1782) );
  OAI222XL U3115 ( .A0(n1054), .A1(n3193), .B0(n4057), .B1(n325), .C0(n4232), 
        .C1(n3954), .Y(n1781) );
  OAI222XL U3116 ( .A0(n1055), .A1(n3193), .B0(n4059), .B1(n325), .C0(n4231), 
        .C1(n3954), .Y(n1780) );
  OAI222XL U3117 ( .A0(n1056), .A1(n3193), .B0(n4062), .B1(n3853), .C0(n4230), 
        .C1(n3954), .Y(n1779) );
  OAI222XL U3118 ( .A0(n1057), .A1(n3193), .B0(n4065), .B1(n3853), .C0(n4229), 
        .C1(n3954), .Y(n1778) );
  OAI222XL U3119 ( .A0(n1058), .A1(n3193), .B0(n4068), .B1(n3853), .C0(n4228), 
        .C1(n3954), .Y(n1777) );
  OAI222XL U3120 ( .A0(n1059), .A1(n3193), .B0(n4071), .B1(n3853), .C0(n4227), 
        .C1(n3954), .Y(n1776) );
  OAI222XL U3121 ( .A0(n1060), .A1(n3193), .B0(n4074), .B1(n3853), .C0(n4226), 
        .C1(n3954), .Y(n1775) );
  OAI222XL U3122 ( .A0(n1061), .A1(n3193), .B0(n4077), .B1(n3853), .C0(n4225), 
        .C1(n3954), .Y(n1774) );
  OAI222XL U3123 ( .A0(n1062), .A1(n3193), .B0(n4080), .B1(n3853), .C0(n4224), 
        .C1(n3954), .Y(n1773) );
  OAI222XL U3124 ( .A0(n1063), .A1(n3193), .B0(n4083), .B1(n3853), .C0(n4223), 
        .C1(n3954), .Y(n1772) );
  OAI222XL U3125 ( .A0(n1064), .A1(n3193), .B0(n4086), .B1(n3853), .C0(n4222), 
        .C1(n3954), .Y(n1771) );
  OAI222XL U3126 ( .A0(n1065), .A1(n3193), .B0(n4089), .B1(n3853), .C0(n4221), 
        .C1(n3954), .Y(n1770) );
  OAI222XL U3127 ( .A0(n1066), .A1(n3193), .B0(n4092), .B1(n3853), .C0(n4220), 
        .C1(n3954), .Y(n1769) );
  OAI222XL U3128 ( .A0(n1067), .A1(n3193), .B0(n4095), .B1(n3853), .C0(n4219), 
        .C1(n3955), .Y(n1768) );
  OAI222XL U3129 ( .A0(n1068), .A1(n3193), .B0(n4098), .B1(n3852), .C0(n4218), 
        .C1(n3955), .Y(n1767) );
  OAI222XL U3130 ( .A0(n1069), .A1(n3193), .B0(n4101), .B1(n3852), .C0(n4217), 
        .C1(n3955), .Y(n1766) );
  OAI222XL U3131 ( .A0(n1070), .A1(n3193), .B0(n4104), .B1(n3852), .C0(n4216), 
        .C1(n3955), .Y(n1765) );
  OAI222XL U3132 ( .A0(n1071), .A1(n3193), .B0(n4107), .B1(n3852), .C0(n4215), 
        .C1(n3955), .Y(n1764) );
  OAI222XL U3133 ( .A0(n1072), .A1(n3193), .B0(n4110), .B1(n3852), .C0(n4214), 
        .C1(n3955), .Y(n1763) );
  OAI222XL U3134 ( .A0(n1073), .A1(n3193), .B0(n4029), .B1(n3852), .C0(n4213), 
        .C1(n3955), .Y(n1762) );
  OAI222XL U3135 ( .A0(n1074), .A1(n3193), .B0(n4031), .B1(n3852), .C0(n4212), 
        .C1(n3955), .Y(n1761) );
  OAI222XL U3136 ( .A0(n1075), .A1(n3193), .B0(n4033), .B1(n3852), .C0(n4211), 
        .C1(n3955), .Y(n1760) );
  OAI222XL U3137 ( .A0(n1076), .A1(n3193), .B0(n4035), .B1(n3852), .C0(n4210), 
        .C1(n3955), .Y(n1759) );
  OAI222XL U3138 ( .A0(n1077), .A1(n3193), .B0(n4037), .B1(n3852), .C0(n4209), 
        .C1(n3955), .Y(n1758) );
  OAI222XL U3139 ( .A0(n1078), .A1(n3193), .B0(n4039), .B1(n3852), .C0(n4208), 
        .C1(n3955), .Y(n1757) );
  OAI222XL U3140 ( .A0(n1079), .A1(n3193), .B0(n4041), .B1(n3852), .C0(n4207), 
        .C1(n3955), .Y(n1756) );
  OAI222XL U3141 ( .A0(n1447), .A1(n4015), .B0(n4044), .B1(n3261), .C0(n4238), 
        .C1(n3862), .Y(n2683) );
  OAI222XL U3142 ( .A0(n1448), .A1(n4015), .B0(n4047), .B1(n3261), .C0(n4237), 
        .C1(n3862), .Y(n2682) );
  OAI222XL U3143 ( .A0(n1449), .A1(n4015), .B0(n4049), .B1(n3261), .C0(n4236), 
        .C1(n3863), .Y(n2681) );
  OAI222XL U3144 ( .A0(n1450), .A1(n4015), .B0(n4051), .B1(n3261), .C0(n4235), 
        .C1(n3863), .Y(n2680) );
  OAI222XL U3145 ( .A0(n1451), .A1(n4015), .B0(n4053), .B1(n3261), .C0(n4234), 
        .C1(n3863), .Y(n2679) );
  OAI222XL U3146 ( .A0(n1452), .A1(n4015), .B0(n4055), .B1(n3261), .C0(n4233), 
        .C1(n3863), .Y(n2678) );
  OAI222XL U3147 ( .A0(n1453), .A1(n4015), .B0(n4057), .B1(n3261), .C0(n4232), 
        .C1(n3863), .Y(n2677) );
  OAI222XL U3148 ( .A0(n1454), .A1(n4015), .B0(n4059), .B1(n3261), .C0(n4231), 
        .C1(n3863), .Y(n2676) );
  OAI222XL U3149 ( .A0(n1455), .A1(n4015), .B0(n4062), .B1(n3261), .C0(n4230), 
        .C1(n3863), .Y(n2675) );
  OAI222XL U3150 ( .A0(n1456), .A1(n4015), .B0(n4065), .B1(n3261), .C0(n4229), 
        .C1(n3863), .Y(n2674) );
  OAI222XL U3151 ( .A0(n1457), .A1(n4015), .B0(n4068), .B1(n3261), .C0(n4228), 
        .C1(n3863), .Y(n2673) );
  OAI222XL U3152 ( .A0(n1458), .A1(n4015), .B0(n4071), .B1(n3261), .C0(n4227), 
        .C1(n3863), .Y(n2672) );
  OAI222XL U3153 ( .A0(n1459), .A1(n4015), .B0(n4074), .B1(n3261), .C0(n4226), 
        .C1(n3863), .Y(n2671) );
  OAI222XL U3154 ( .A0(n1460), .A1(n4015), .B0(n4077), .B1(n3261), .C0(n4225), 
        .C1(n3863), .Y(n2670) );
  OAI222XL U3155 ( .A0(n1461), .A1(n4015), .B0(n4080), .B1(n3261), .C0(n4224), 
        .C1(n3863), .Y(n2669) );
  OAI222XL U3156 ( .A0(n1462), .A1(n4015), .B0(n4083), .B1(n3261), .C0(n4223), 
        .C1(n3863), .Y(n2668) );
  OAI222XL U3157 ( .A0(n1463), .A1(n4015), .B0(n4086), .B1(n3261), .C0(n4222), 
        .C1(n3863), .Y(n2667) );
  OAI222XL U3158 ( .A0(n1464), .A1(n4015), .B0(n4089), .B1(n3261), .C0(n4221), 
        .C1(n3863), .Y(n2666) );
  OAI222XL U3159 ( .A0(n1465), .A1(n4015), .B0(n4092), .B1(n3261), .C0(n4220), 
        .C1(n3864), .Y(n2665) );
  OAI222XL U3160 ( .A0(n1466), .A1(n4015), .B0(n4095), .B1(n3261), .C0(n4219), 
        .C1(n3864), .Y(n2664) );
  OAI222XL U3161 ( .A0(n1467), .A1(n4015), .B0(n4098), .B1(n3261), .C0(n4218), 
        .C1(n3864), .Y(n2663) );
  OAI222XL U3162 ( .A0(n1468), .A1(n4015), .B0(n4101), .B1(n3261), .C0(n4217), 
        .C1(n3864), .Y(n2662) );
  OAI222XL U3163 ( .A0(n1469), .A1(n4015), .B0(n4104), .B1(n3261), .C0(n4216), 
        .C1(n3864), .Y(n2661) );
  OAI222XL U3164 ( .A0(n1470), .A1(n4015), .B0(n4107), .B1(n3261), .C0(n4215), 
        .C1(n3864), .Y(n2660) );
  OAI222XL U3165 ( .A0(n1471), .A1(n4015), .B0(n4110), .B1(n3261), .C0(n4214), 
        .C1(n3864), .Y(n2659) );
  OAI222XL U3166 ( .A0(n1472), .A1(n4015), .B0(n4028), .B1(n3261), .C0(n4213), 
        .C1(n3864), .Y(n2658) );
  OAI222XL U3167 ( .A0(n1473), .A1(n4015), .B0(n4030), .B1(n3261), .C0(n4212), 
        .C1(n3864), .Y(n2657) );
  OAI222XL U3168 ( .A0(n1474), .A1(n4015), .B0(n4032), .B1(n3261), .C0(n4211), 
        .C1(n3864), .Y(n2656) );
  OAI222XL U3169 ( .A0(n1475), .A1(n4015), .B0(n4034), .B1(n3261), .C0(n4210), 
        .C1(n3864), .Y(n2655) );
  OAI222XL U3170 ( .A0(n1476), .A1(n4015), .B0(n4036), .B1(n3261), .C0(n4209), 
        .C1(n3864), .Y(n2654) );
  OAI222XL U3171 ( .A0(n1477), .A1(n4015), .B0(n4038), .B1(n3261), .C0(n4208), 
        .C1(n3864), .Y(n2653) );
  OAI222XL U3172 ( .A0(n1478), .A1(n4015), .B0(n4040), .B1(n3261), .C0(n4207), 
        .C1(n3864), .Y(n2652) );
  OAI222XL U3173 ( .A0(n1575), .A1(n4026), .B0(n4044), .B1(n3185), .C0(n3876), 
        .C1(n4238), .Y(n2555) );
  OAI222XL U3174 ( .A0(n1576), .A1(n4026), .B0(n4047), .B1(n3185), .C0(n3876), 
        .C1(n4237), .Y(n2554) );
  OAI222XL U3175 ( .A0(n1577), .A1(n4026), .B0(n4049), .B1(n3185), .C0(n3876), 
        .C1(n4236), .Y(n2553) );
  OAI222XL U3176 ( .A0(n1578), .A1(n4026), .B0(n4051), .B1(n3185), .C0(n3876), 
        .C1(n4235), .Y(n2552) );
  OAI222XL U3177 ( .A0(n1579), .A1(n4026), .B0(n4053), .B1(n3185), .C0(n3877), 
        .C1(n4234), .Y(n2551) );
  OAI222XL U3178 ( .A0(n1580), .A1(n4026), .B0(n4055), .B1(n3185), .C0(n3877), 
        .C1(n4233), .Y(n2550) );
  OAI222XL U3179 ( .A0(n1581), .A1(n4026), .B0(n4057), .B1(n3185), .C0(n3877), 
        .C1(n4232), .Y(n2549) );
  OAI222XL U3180 ( .A0(n1582), .A1(n4026), .B0(n4059), .B1(n3185), .C0(n3877), 
        .C1(n4231), .Y(n2548) );
  OAI222XL U3181 ( .A0(n1583), .A1(n4026), .B0(n4062), .B1(n3185), .C0(n3877), 
        .C1(n4230), .Y(n2547) );
  OAI222XL U3182 ( .A0(n1584), .A1(n4026), .B0(n4065), .B1(n3185), .C0(n3877), 
        .C1(n4229), .Y(n2546) );
  OAI222XL U3183 ( .A0(n1585), .A1(n4026), .B0(n4068), .B1(n3185), .C0(n3877), 
        .C1(n4228), .Y(n2545) );
  OAI222XL U3184 ( .A0(n1586), .A1(n4026), .B0(n4071), .B1(n3185), .C0(n3877), 
        .C1(n4227), .Y(n2544) );
  OAI222XL U3185 ( .A0(n1587), .A1(n4026), .B0(n4074), .B1(n3185), .C0(n3877), 
        .C1(n4226), .Y(n2543) );
  OAI222XL U3186 ( .A0(n1588), .A1(n4026), .B0(n4077), .B1(n3185), .C0(n3877), 
        .C1(n4225), .Y(n2542) );
  OAI222XL U3187 ( .A0(n1589), .A1(n4026), .B0(n4080), .B1(n3185), .C0(n3877), 
        .C1(n4224), .Y(n2541) );
  OAI222XL U3188 ( .A0(n1590), .A1(n4026), .B0(n4083), .B1(n3185), .C0(n3877), 
        .C1(n4223), .Y(n2540) );
  OAI222XL U3189 ( .A0(n1591), .A1(n4026), .B0(n4086), .B1(n3185), .C0(n3877), 
        .C1(n4222), .Y(n2539) );
  OAI222XL U3190 ( .A0(n1592), .A1(n4026), .B0(n4089), .B1(n3185), .C0(n3877), 
        .C1(n4221), .Y(n2538) );
  OAI222XL U3191 ( .A0(n1593), .A1(n4026), .B0(n4092), .B1(n3185), .C0(n3877), 
        .C1(n4220), .Y(n2537) );
  OAI222XL U3192 ( .A0(n1594), .A1(n4026), .B0(n4095), .B1(n3185), .C0(n3877), 
        .C1(n4219), .Y(n2536) );
  OAI222XL U3193 ( .A0(n1595), .A1(n4026), .B0(n4098), .B1(n3185), .C0(n3878), 
        .C1(n4218), .Y(n2535) );
  OAI222XL U3194 ( .A0(n1596), .A1(n4026), .B0(n4101), .B1(n3185), .C0(n3878), 
        .C1(n4217), .Y(n2534) );
  OAI222XL U3195 ( .A0(n1597), .A1(n4026), .B0(n4104), .B1(n3185), .C0(n3878), 
        .C1(n4216), .Y(n2533) );
  OAI222XL U3196 ( .A0(n1598), .A1(n4026), .B0(n4107), .B1(n3185), .C0(n3878), 
        .C1(n4215), .Y(n2532) );
  OAI222XL U3197 ( .A0(n1599), .A1(n4026), .B0(n4110), .B1(n3185), .C0(n3878), 
        .C1(n4214), .Y(n2531) );
  OAI222XL U3198 ( .A0(n1600), .A1(n4026), .B0(n4029), .B1(n3185), .C0(n3878), 
        .C1(n4213), .Y(n2530) );
  OAI222XL U3199 ( .A0(n1601), .A1(n4026), .B0(n4031), .B1(n3185), .C0(n3878), 
        .C1(n4212), .Y(n2529) );
  OAI222XL U3200 ( .A0(n1602), .A1(n4026), .B0(n4033), .B1(n3185), .C0(n3878), 
        .C1(n4211), .Y(n2528) );
  OAI222XL U3201 ( .A0(n1603), .A1(n4026), .B0(n4035), .B1(n3185), .C0(n3878), 
        .C1(n4210), .Y(n2527) );
  OAI222XL U3202 ( .A0(n1604), .A1(n4026), .B0(n4037), .B1(n3185), .C0(n3878), 
        .C1(n4209), .Y(n2526) );
  OAI222XL U3203 ( .A0(n1605), .A1(n4026), .B0(n4039), .B1(n3185), .C0(n3878), 
        .C1(n4208), .Y(n2525) );
  OAI222XL U3204 ( .A0(n1606), .A1(n4026), .B0(n4041), .B1(n3185), .C0(n3878), 
        .C1(n4207), .Y(n2524) );
  OAI222XL U3205 ( .A0(n440), .A1(n3201), .B0(n4043), .B1(n3815), .C0(n3885), 
        .C1(n4206), .Y(n2395) );
  OAI222XL U3206 ( .A0(n441), .A1(n3201), .B0(n4046), .B1(n3814), .C0(n3886), 
        .C1(n4205), .Y(n2394) );
  OAI222XL U3207 ( .A0(n442), .A1(n3201), .B0(n3203), .B1(n365), .C0(n3885), 
        .C1(n4204), .Y(n2393) );
  OAI222XL U3208 ( .A0(n443), .A1(n3201), .B0(n3204), .B1(n365), .C0(n3885), 
        .C1(n4203), .Y(n2392) );
  OAI222XL U3209 ( .A0(n444), .A1(n3201), .B0(n3210), .B1(n365), .C0(n3886), 
        .C1(n4202), .Y(n2391) );
  OAI222XL U3210 ( .A0(n445), .A1(n3201), .B0(n3211), .B1(n365), .C0(n3885), 
        .C1(n4201), .Y(n2390) );
  OAI222XL U3211 ( .A0(n446), .A1(n3201), .B0(n3212), .B1(n365), .C0(n3885), 
        .C1(n4200), .Y(n2389) );
  OAI222XL U3212 ( .A0(n447), .A1(n3201), .B0(n3213), .B1(n365), .C0(n3886), 
        .C1(n4199), .Y(n2388) );
  OAI222XL U3213 ( .A0(n448), .A1(n3201), .B0(n4061), .B1(n3815), .C0(n3885), 
        .C1(n4198), .Y(n2387) );
  OAI222XL U3214 ( .A0(n449), .A1(n3201), .B0(n4064), .B1(n3815), .C0(n3886), 
        .C1(n4197), .Y(n2386) );
  OAI222XL U3215 ( .A0(n450), .A1(n3201), .B0(n4067), .B1(n3815), .C0(n3886), 
        .C1(n4196), .Y(n2385) );
  OAI222XL U3216 ( .A0(n451), .A1(n3201), .B0(n4070), .B1(n3815), .C0(n3886), 
        .C1(n4195), .Y(n2384) );
  OAI222XL U3217 ( .A0(n452), .A1(n3201), .B0(n4073), .B1(n3815), .C0(n3886), 
        .C1(n4194), .Y(n2383) );
  OAI222XL U3218 ( .A0(n453), .A1(n3201), .B0(n4076), .B1(n3815), .C0(n3887), 
        .C1(n4193), .Y(n2382) );
  OAI222XL U3219 ( .A0(n454), .A1(n3201), .B0(n4079), .B1(n3815), .C0(n3887), 
        .C1(n4192), .Y(n2381) );
  OAI222XL U3220 ( .A0(n455), .A1(n3201), .B0(n4082), .B1(n3815), .C0(n3887), 
        .C1(n4191), .Y(n2380) );
  OAI222XL U3221 ( .A0(n456), .A1(n3201), .B0(n4085), .B1(n3815), .C0(n3887), 
        .C1(n4190), .Y(n2379) );
  OAI222XL U3222 ( .A0(n457), .A1(n3201), .B0(n4088), .B1(n3815), .C0(n3887), 
        .C1(n4189), .Y(n2378) );
  OAI222XL U3223 ( .A0(n458), .A1(n3201), .B0(n4091), .B1(n3815), .C0(n3887), 
        .C1(n4188), .Y(n2377) );
  OAI222XL U3224 ( .A0(n459), .A1(n3201), .B0(n4094), .B1(n3815), .C0(n3887), 
        .C1(n4187), .Y(n2376) );
  OAI222XL U3225 ( .A0(n460), .A1(n3201), .B0(n4097), .B1(n3814), .C0(n3887), 
        .C1(n4186), .Y(n2375) );
  OAI222XL U3226 ( .A0(n461), .A1(n3201), .B0(n4100), .B1(n3814), .C0(n3887), 
        .C1(n4185), .Y(n2374) );
  OAI222XL U3227 ( .A0(n462), .A1(n3201), .B0(n4103), .B1(n3814), .C0(n3887), 
        .C1(n4184), .Y(n2373) );
  OAI222XL U3228 ( .A0(n463), .A1(n3201), .B0(n4106), .B1(n3814), .C0(n3887), 
        .C1(n4183), .Y(n2372) );
  OAI222XL U3229 ( .A0(n464), .A1(n3201), .B0(n3209), .B1(n3814), .C0(n3887), 
        .C1(n4182), .Y(n2371) );
  OAI222XL U3230 ( .A0(n465), .A1(n3201), .B0(n4028), .B1(n3814), .C0(n3887), 
        .C1(n4181), .Y(n2370) );
  OAI222XL U3231 ( .A0(n466), .A1(n3201), .B0(n4030), .B1(n3814), .C0(n3887), 
        .C1(n4180), .Y(n2369) );
  OAI222XL U3232 ( .A0(n467), .A1(n3201), .B0(n4032), .B1(n3814), .C0(n3887), 
        .C1(n4179), .Y(n2368) );
  OAI222XL U3233 ( .A0(n468), .A1(n3201), .B0(n4034), .B1(n3814), .C0(n3888), 
        .C1(n4178), .Y(n2367) );
  OAI222XL U3234 ( .A0(n469), .A1(n3201), .B0(n4036), .B1(n3814), .C0(n3888), 
        .C1(n4177), .Y(n2366) );
  OAI222XL U3235 ( .A0(n470), .A1(n3201), .B0(n4038), .B1(n3814), .C0(n3888), 
        .C1(n4176), .Y(n2365) );
  OAI222XL U3236 ( .A0(n471), .A1(n3201), .B0(n4040), .B1(n3814), .C0(n3888), 
        .C1(n4175), .Y(n2364) );
  OAI222XL U3237 ( .A0(n568), .A1(n3187), .B0(n4043), .B1(n3823), .C0(n4206), 
        .C1(n3903), .Y(n2267) );
  OAI222XL U3238 ( .A0(n569), .A1(n3187), .B0(n4046), .B1(n3822), .C0(n4205), 
        .C1(n3903), .Y(n2266) );
  OAI222XL U3239 ( .A0(n570), .A1(n3187), .B0(n4050), .B1(n355), .C0(n4204), 
        .C1(n3903), .Y(n2265) );
  OAI222XL U3240 ( .A0(n571), .A1(n3187), .B0(n4052), .B1(n355), .C0(n4203), 
        .C1(n3904), .Y(n2264) );
  OAI222XL U3241 ( .A0(n572), .A1(n3187), .B0(n4054), .B1(n355), .C0(n4202), 
        .C1(n3904), .Y(n2263) );
  OAI222XL U3242 ( .A0(n573), .A1(n3187), .B0(n4056), .B1(n355), .C0(n4201), 
        .C1(n3904), .Y(n2262) );
  OAI222XL U3243 ( .A0(n574), .A1(n3187), .B0(n4058), .B1(n355), .C0(n4200), 
        .C1(n3904), .Y(n2261) );
  OAI222XL U3244 ( .A0(n575), .A1(n3187), .B0(n4060), .B1(n355), .C0(n4199), 
        .C1(n3904), .Y(n2260) );
  OAI222XL U3245 ( .A0(n576), .A1(n3187), .B0(n4061), .B1(n3823), .C0(n4198), 
        .C1(n3904), .Y(n2259) );
  OAI222XL U3246 ( .A0(n577), .A1(n3187), .B0(n4064), .B1(n3823), .C0(n4197), 
        .C1(n3904), .Y(n2258) );
  OAI222XL U3247 ( .A0(n578), .A1(n3187), .B0(n4067), .B1(n3823), .C0(n4196), 
        .C1(n3904), .Y(n2257) );
  OAI222XL U3248 ( .A0(n579), .A1(n3187), .B0(n4070), .B1(n3823), .C0(n4195), 
        .C1(n3904), .Y(n2256) );
  OAI222XL U3249 ( .A0(n580), .A1(n3187), .B0(n4073), .B1(n3823), .C0(n4194), 
        .C1(n3904), .Y(n2255) );
  OAI222XL U3250 ( .A0(n581), .A1(n3187), .B0(n4076), .B1(n3823), .C0(n4193), 
        .C1(n3904), .Y(n2254) );
  OAI222XL U3251 ( .A0(n582), .A1(n3187), .B0(n4079), .B1(n3823), .C0(n4192), 
        .C1(n3904), .Y(n2253) );
  OAI222XL U3252 ( .A0(n583), .A1(n3187), .B0(n4082), .B1(n3823), .C0(n4191), 
        .C1(n3904), .Y(n2252) );
  OAI222XL U3253 ( .A0(n584), .A1(n3187), .B0(n4085), .B1(n3823), .C0(n4190), 
        .C1(n3904), .Y(n2251) );
  OAI222XL U3254 ( .A0(n585), .A1(n3187), .B0(n4088), .B1(n3823), .C0(n4189), 
        .C1(n3904), .Y(n2250) );
  OAI222XL U3255 ( .A0(n586), .A1(n3187), .B0(n4091), .B1(n3823), .C0(n4188), 
        .C1(n3904), .Y(n2249) );
  OAI222XL U3256 ( .A0(n587), .A1(n3187), .B0(n4094), .B1(n3823), .C0(n4187), 
        .C1(n3897), .Y(n2248) );
  OAI222XL U3257 ( .A0(n588), .A1(n3187), .B0(n4097), .B1(n3822), .C0(n4186), 
        .C1(n3904), .Y(n2247) );
  OAI222XL U3258 ( .A0(n589), .A1(n3187), .B0(n4100), .B1(n3822), .C0(n4185), 
        .C1(n3897), .Y(n2246) );
  OAI222XL U3259 ( .A0(n590), .A1(n3187), .B0(n4103), .B1(n3822), .C0(n4184), 
        .C1(n3901), .Y(n2245) );
  OAI222XL U3260 ( .A0(n591), .A1(n3187), .B0(n4106), .B1(n3822), .C0(n4183), 
        .C1(n3903), .Y(n2244) );
  OAI222XL U3261 ( .A0(n592), .A1(n3187), .B0(n3209), .B1(n3822), .C0(n4182), 
        .C1(n3897), .Y(n2243) );
  OAI222XL U3262 ( .A0(n593), .A1(n3187), .B0(n4028), .B1(n3822), .C0(n4181), 
        .C1(n3897), .Y(n2242) );
  OAI222XL U3263 ( .A0(n594), .A1(n3187), .B0(n4030), .B1(n3822), .C0(n4180), 
        .C1(n3899), .Y(n2241) );
  OAI222XL U3264 ( .A0(n595), .A1(n3187), .B0(n4032), .B1(n3822), .C0(n4179), 
        .C1(n3903), .Y(n2240) );
  OAI222XL U3265 ( .A0(n596), .A1(n3187), .B0(n4034), .B1(n3822), .C0(n4178), 
        .C1(n3897), .Y(n2239) );
  OAI222XL U3266 ( .A0(n597), .A1(n3187), .B0(n4036), .B1(n3822), .C0(n4177), 
        .C1(n3897), .Y(n2238) );
  OAI222XL U3267 ( .A0(n598), .A1(n3187), .B0(n4038), .B1(n3822), .C0(n4176), 
        .C1(n3897), .Y(n2237) );
  OAI222XL U3268 ( .A0(n599), .A1(n3187), .B0(n4040), .B1(n3822), .C0(n4175), 
        .C1(n3899), .Y(n2236) );
  OAI222XL U3269 ( .A0(n696), .A1(n3186), .B0(n4045), .B1(n3831), .C0(n4206), 
        .C1(n3916), .Y(n2139) );
  OAI222XL U3270 ( .A0(n697), .A1(n3186), .B0(n4048), .B1(n3830), .C0(n4205), 
        .C1(n3916), .Y(n2138) );
  OAI222XL U3271 ( .A0(n698), .A1(n3186), .B0(n4050), .B1(n347), .C0(n4204), 
        .C1(n3916), .Y(n2137) );
  OAI222XL U3272 ( .A0(n699), .A1(n3186), .B0(n4052), .B1(n347), .C0(n4203), 
        .C1(n3917), .Y(n2136) );
  OAI222XL U3273 ( .A0(n700), .A1(n3186), .B0(n4054), .B1(n347), .C0(n4202), 
        .C1(n3917), .Y(n2135) );
  OAI222XL U3274 ( .A0(n701), .A1(n3186), .B0(n4056), .B1(n347), .C0(n4201), 
        .C1(n3917), .Y(n2134) );
  OAI222XL U3275 ( .A0(n702), .A1(n3186), .B0(n4058), .B1(n347), .C0(n4200), 
        .C1(n3917), .Y(n2133) );
  OAI222XL U3276 ( .A0(n703), .A1(n3186), .B0(n4060), .B1(n347), .C0(n4199), 
        .C1(n3917), .Y(n2132) );
  OAI222XL U3277 ( .A0(n704), .A1(n3186), .B0(n4063), .B1(n3831), .C0(n4198), 
        .C1(n3917), .Y(n2131) );
  OAI222XL U3278 ( .A0(n705), .A1(n3186), .B0(n4066), .B1(n3831), .C0(n4197), 
        .C1(n3917), .Y(n2130) );
  OAI222XL U3279 ( .A0(n706), .A1(n3186), .B0(n4069), .B1(n3831), .C0(n4196), 
        .C1(n3917), .Y(n2129) );
  OAI222XL U3280 ( .A0(n707), .A1(n3186), .B0(n4072), .B1(n3831), .C0(n4195), 
        .C1(n3917), .Y(n2128) );
  OAI222XL U3281 ( .A0(n708), .A1(n3186), .B0(n4075), .B1(n3831), .C0(n4194), 
        .C1(n3917), .Y(n2127) );
  OAI222XL U3282 ( .A0(n709), .A1(n3186), .B0(n4078), .B1(n3831), .C0(n4193), 
        .C1(n3917), .Y(n2126) );
  OAI222XL U3283 ( .A0(n710), .A1(n3186), .B0(n4081), .B1(n3831), .C0(n4192), 
        .C1(n3917), .Y(n2125) );
  OAI222XL U3284 ( .A0(n711), .A1(n3186), .B0(n4084), .B1(n3831), .C0(n4191), 
        .C1(n3917), .Y(n2124) );
  OAI222XL U3285 ( .A0(n712), .A1(n3186), .B0(n4087), .B1(n3831), .C0(n4190), 
        .C1(n3917), .Y(n2123) );
  OAI222XL U3286 ( .A0(n713), .A1(n3186), .B0(n4090), .B1(n3831), .C0(n4189), 
        .C1(n3917), .Y(n2122) );
  OAI222XL U3287 ( .A0(n714), .A1(n3186), .B0(n4093), .B1(n3831), .C0(n4188), 
        .C1(n3917), .Y(n2121) );
  OAI222XL U3288 ( .A0(n715), .A1(n3186), .B0(n4096), .B1(n3831), .C0(n4187), 
        .C1(n3910), .Y(n2120) );
  OAI222XL U3289 ( .A0(n716), .A1(n3186), .B0(n4099), .B1(n3830), .C0(n4186), 
        .C1(n3917), .Y(n2119) );
  OAI222XL U3290 ( .A0(n717), .A1(n3186), .B0(n4102), .B1(n3830), .C0(n4185), 
        .C1(n3910), .Y(n2118) );
  OAI222XL U3291 ( .A0(n718), .A1(n3186), .B0(n4105), .B1(n3830), .C0(n4184), 
        .C1(n3917), .Y(n2117) );
  OAI222XL U3292 ( .A0(n719), .A1(n3186), .B0(n4108), .B1(n3830), .C0(n4183), 
        .C1(n3916), .Y(n2116) );
  OAI222XL U3293 ( .A0(n720), .A1(n3186), .B0(n4111), .B1(n3830), .C0(n4182), 
        .C1(n3910), .Y(n2115) );
  OAI222XL U3294 ( .A0(n721), .A1(n3186), .B0(n4028), .B1(n3830), .C0(n4181), 
        .C1(n3910), .Y(n2114) );
  OAI222XL U3295 ( .A0(n722), .A1(n3186), .B0(n4030), .B1(n3830), .C0(n4180), 
        .C1(n3912), .Y(n2113) );
  OAI222XL U3296 ( .A0(n723), .A1(n3186), .B0(n4032), .B1(n3830), .C0(n4179), 
        .C1(n3916), .Y(n2112) );
  OAI222XL U3297 ( .A0(n724), .A1(n3186), .B0(n4034), .B1(n3830), .C0(n4178), 
        .C1(n3910), .Y(n2111) );
  OAI222XL U3298 ( .A0(n725), .A1(n3186), .B0(n4036), .B1(n3830), .C0(n4177), 
        .C1(n3910), .Y(n2110) );
  OAI222XL U3299 ( .A0(n726), .A1(n3186), .B0(n4038), .B1(n3830), .C0(n4176), 
        .C1(n3910), .Y(n2109) );
  OAI222XL U3300 ( .A0(n727), .A1(n3186), .B0(n4040), .B1(n3830), .C0(n4175), 
        .C1(n3912), .Y(n2108) );
  OAI222XL U3301 ( .A0(n824), .A1(n3190), .B0(n4045), .B1(n3839), .C0(n4206), 
        .C1(n3929), .Y(n2011) );
  OAI222XL U3302 ( .A0(n825), .A1(n3190), .B0(n4048), .B1(n3838), .C0(n4205), 
        .C1(n3929), .Y(n2010) );
  OAI222XL U3303 ( .A0(n826), .A1(n3190), .B0(n4050), .B1(n339), .C0(n4204), 
        .C1(n3929), .Y(n2009) );
  OAI222XL U3304 ( .A0(n827), .A1(n3190), .B0(n4052), .B1(n339), .C0(n4203), 
        .C1(n3930), .Y(n2008) );
  OAI222XL U3305 ( .A0(n828), .A1(n3190), .B0(n4054), .B1(n339), .C0(n4202), 
        .C1(n3930), .Y(n2007) );
  OAI222XL U3306 ( .A0(n829), .A1(n3190), .B0(n4056), .B1(n339), .C0(n4201), 
        .C1(n3930), .Y(n2006) );
  OAI222XL U3307 ( .A0(n830), .A1(n3190), .B0(n4058), .B1(n339), .C0(n4200), 
        .C1(n3930), .Y(n2005) );
  OAI222XL U3308 ( .A0(n831), .A1(n3190), .B0(n4060), .B1(n339), .C0(n4199), 
        .C1(n3930), .Y(n2004) );
  OAI222XL U3309 ( .A0(n832), .A1(n3190), .B0(n4063), .B1(n3839), .C0(n4198), 
        .C1(n3930), .Y(n2003) );
  OAI222XL U3310 ( .A0(n833), .A1(n3190), .B0(n4066), .B1(n3839), .C0(n4197), 
        .C1(n3930), .Y(n2002) );
  OAI222XL U3311 ( .A0(n834), .A1(n3190), .B0(n4069), .B1(n3839), .C0(n4196), 
        .C1(n3930), .Y(n2001) );
  OAI222XL U3312 ( .A0(n835), .A1(n3190), .B0(n4072), .B1(n3839), .C0(n4195), 
        .C1(n3930), .Y(n2000) );
  OAI222XL U3313 ( .A0(n836), .A1(n3190), .B0(n4075), .B1(n3839), .C0(n4194), 
        .C1(n3930), .Y(n1999) );
  OAI222XL U3314 ( .A0(n837), .A1(n3190), .B0(n4078), .B1(n3839), .C0(n4193), 
        .C1(n3930), .Y(n1998) );
  OAI222XL U3315 ( .A0(n838), .A1(n3190), .B0(n4081), .B1(n3839), .C0(n4192), 
        .C1(n3930), .Y(n1997) );
  OAI222XL U3316 ( .A0(n839), .A1(n3190), .B0(n4084), .B1(n3839), .C0(n4191), 
        .C1(n3930), .Y(n1996) );
  OAI222XL U3317 ( .A0(n840), .A1(n3190), .B0(n4087), .B1(n3839), .C0(n4190), 
        .C1(n3930), .Y(n1995) );
  OAI222XL U3318 ( .A0(n841), .A1(n3190), .B0(n4090), .B1(n3839), .C0(n4189), 
        .C1(n3930), .Y(n1994) );
  OAI222XL U3319 ( .A0(n842), .A1(n3190), .B0(n4093), .B1(n3839), .C0(n4188), 
        .C1(n3930), .Y(n1993) );
  OAI222XL U3320 ( .A0(n843), .A1(n3190), .B0(n4096), .B1(n3839), .C0(n4187), 
        .C1(n3923), .Y(n1992) );
  OAI222XL U3321 ( .A0(n844), .A1(n3190), .B0(n4099), .B1(n3838), .C0(n4186), 
        .C1(n3930), .Y(n1991) );
  OAI222XL U3322 ( .A0(n845), .A1(n3190), .B0(n4102), .B1(n3838), .C0(n4185), 
        .C1(n3923), .Y(n1990) );
  OAI222XL U3323 ( .A0(n846), .A1(n3190), .B0(n4105), .B1(n3838), .C0(n4184), 
        .C1(n3930), .Y(n1989) );
  OAI222XL U3324 ( .A0(n847), .A1(n3190), .B0(n4108), .B1(n3838), .C0(n4183), 
        .C1(n3929), .Y(n1988) );
  OAI222XL U3325 ( .A0(n848), .A1(n3190), .B0(n4111), .B1(n3838), .C0(n4182), 
        .C1(n3923), .Y(n1987) );
  OAI222XL U3326 ( .A0(n849), .A1(n3190), .B0(n4029), .B1(n3838), .C0(n4181), 
        .C1(n3929), .Y(n1986) );
  OAI222XL U3327 ( .A0(n850), .A1(n3190), .B0(n4031), .B1(n3838), .C0(n4180), 
        .C1(n3923), .Y(n1985) );
  OAI222XL U3328 ( .A0(n851), .A1(n3190), .B0(n4033), .B1(n3838), .C0(n4179), 
        .C1(n3925), .Y(n1984) );
  OAI222XL U3329 ( .A0(n852), .A1(n3190), .B0(n4035), .B1(n3838), .C0(n4178), 
        .C1(n3923), .Y(n1983) );
  OAI222XL U3330 ( .A0(n853), .A1(n3190), .B0(n4037), .B1(n3838), .C0(n4177), 
        .C1(n3923), .Y(n1982) );
  OAI222XL U3331 ( .A0(n854), .A1(n3190), .B0(n4039), .B1(n3838), .C0(n4176), 
        .C1(n3923), .Y(n1981) );
  OAI222XL U3332 ( .A0(n855), .A1(n3190), .B0(n4041), .B1(n3838), .C0(n4175), 
        .C1(n3925), .Y(n1980) );
  OAI222XL U3333 ( .A0(n952), .A1(n3189), .B0(n4045), .B1(n3847), .C0(n4206), 
        .C1(n3942), .Y(n1883) );
  OAI222XL U3334 ( .A0(n953), .A1(n3189), .B0(n4048), .B1(n3846), .C0(n4205), 
        .C1(n3942), .Y(n1882) );
  OAI222XL U3335 ( .A0(n954), .A1(n3189), .B0(n4050), .B1(n331), .C0(n4204), 
        .C1(n3942), .Y(n1881) );
  OAI222XL U3336 ( .A0(n955), .A1(n3189), .B0(n4052), .B1(n331), .C0(n4203), 
        .C1(n3943), .Y(n1880) );
  OAI222XL U3337 ( .A0(n956), .A1(n3189), .B0(n4054), .B1(n331), .C0(n4202), 
        .C1(n3943), .Y(n1879) );
  OAI222XL U3338 ( .A0(n957), .A1(n3189), .B0(n4056), .B1(n331), .C0(n4201), 
        .C1(n3943), .Y(n1878) );
  OAI222XL U3339 ( .A0(n958), .A1(n3189), .B0(n4058), .B1(n331), .C0(n4200), 
        .C1(n3943), .Y(n1877) );
  OAI222XL U3340 ( .A0(n959), .A1(n3189), .B0(n4060), .B1(n331), .C0(n4199), 
        .C1(n3943), .Y(n1876) );
  OAI222XL U3341 ( .A0(n960), .A1(n3189), .B0(n4063), .B1(n3847), .C0(n4198), 
        .C1(n3943), .Y(n1875) );
  OAI222XL U3342 ( .A0(n961), .A1(n3189), .B0(n4066), .B1(n3847), .C0(n4197), 
        .C1(n3943), .Y(n1874) );
  OAI222XL U3343 ( .A0(n962), .A1(n3189), .B0(n4069), .B1(n3847), .C0(n4196), 
        .C1(n3943), .Y(n1873) );
  OAI222XL U3344 ( .A0(n963), .A1(n3189), .B0(n4072), .B1(n3847), .C0(n4195), 
        .C1(n3943), .Y(n1872) );
  OAI222XL U3345 ( .A0(n964), .A1(n3189), .B0(n4075), .B1(n3847), .C0(n4194), 
        .C1(n3943), .Y(n1871) );
  OAI222XL U3346 ( .A0(n965), .A1(n3189), .B0(n4078), .B1(n3847), .C0(n4193), 
        .C1(n3943), .Y(n1870) );
  OAI222XL U3347 ( .A0(n966), .A1(n3189), .B0(n4081), .B1(n3847), .C0(n4192), 
        .C1(n3943), .Y(n1869) );
  OAI222XL U3348 ( .A0(n967), .A1(n3189), .B0(n4084), .B1(n3847), .C0(n4191), 
        .C1(n3943), .Y(n1868) );
  OAI222XL U3349 ( .A0(n968), .A1(n3189), .B0(n4087), .B1(n3847), .C0(n4190), 
        .C1(n3943), .Y(n1867) );
  OAI222XL U3350 ( .A0(n969), .A1(n3189), .B0(n4090), .B1(n3847), .C0(n4189), 
        .C1(n3943), .Y(n1866) );
  OAI222XL U3351 ( .A0(n970), .A1(n3189), .B0(n4093), .B1(n3847), .C0(n4188), 
        .C1(n3943), .Y(n1865) );
  OAI222XL U3352 ( .A0(n971), .A1(n3189), .B0(n4096), .B1(n3847), .C0(n4187), 
        .C1(n3936), .Y(n1864) );
  OAI222XL U3353 ( .A0(n972), .A1(n3189), .B0(n4099), .B1(n3846), .C0(n4186), 
        .C1(n3943), .Y(n1863) );
  OAI222XL U3354 ( .A0(n973), .A1(n3189), .B0(n4102), .B1(n3846), .C0(n4185), 
        .C1(n3936), .Y(n1862) );
  OAI222XL U3355 ( .A0(n974), .A1(n3189), .B0(n4105), .B1(n3846), .C0(n4184), 
        .C1(n3943), .Y(n1861) );
  OAI222XL U3356 ( .A0(n975), .A1(n3189), .B0(n4108), .B1(n3846), .C0(n4183), 
        .C1(n3942), .Y(n1860) );
  OAI222XL U3357 ( .A0(n976), .A1(n3189), .B0(n4111), .B1(n3846), .C0(n4182), 
        .C1(n3936), .Y(n1859) );
  OAI222XL U3358 ( .A0(n977), .A1(n3189), .B0(n4029), .B1(n3846), .C0(n4181), 
        .C1(n3938), .Y(n1858) );
  OAI222XL U3359 ( .A0(n978), .A1(n3189), .B0(n4031), .B1(n3846), .C0(n4180), 
        .C1(n3936), .Y(n1857) );
  OAI222XL U3360 ( .A0(n979), .A1(n3189), .B0(n4033), .B1(n3846), .C0(n4179), 
        .C1(n3942), .Y(n1856) );
  OAI222XL U3361 ( .A0(n980), .A1(n3189), .B0(n4035), .B1(n3846), .C0(n4178), 
        .C1(n3936), .Y(n1855) );
  OAI222XL U3362 ( .A0(n981), .A1(n3189), .B0(n4037), .B1(n3846), .C0(n4177), 
        .C1(n3936), .Y(n1854) );
  OAI222XL U3363 ( .A0(n982), .A1(n3189), .B0(n4039), .B1(n3846), .C0(n4176), 
        .C1(n3936), .Y(n1853) );
  OAI222XL U3364 ( .A0(n983), .A1(n3189), .B0(n4041), .B1(n3846), .C0(n4175), 
        .C1(n3938), .Y(n1852) );
  OAI222XL U3365 ( .A0(n1080), .A1(n3188), .B0(n4044), .B1(n3855), .C0(n4206), 
        .C1(n3955), .Y(n1755) );
  OAI222XL U3366 ( .A0(n1081), .A1(n3188), .B0(n4047), .B1(n3854), .C0(n4205), 
        .C1(n3955), .Y(n1754) );
  OAI222XL U3367 ( .A0(n1082), .A1(n3188), .B0(n4049), .B1(n323), .C0(n4204), 
        .C1(n3955), .Y(n1753) );
  OAI222XL U3368 ( .A0(n1083), .A1(n3188), .B0(n4051), .B1(n323), .C0(n4203), 
        .C1(n3956), .Y(n1752) );
  OAI222XL U3369 ( .A0(n1084), .A1(n3188), .B0(n4053), .B1(n323), .C0(n4202), 
        .C1(n3956), .Y(n1751) );
  OAI222XL U3370 ( .A0(n1085), .A1(n3188), .B0(n4055), .B1(n323), .C0(n4201), 
        .C1(n3956), .Y(n1750) );
  OAI222XL U3371 ( .A0(n1086), .A1(n3188), .B0(n4057), .B1(n323), .C0(n4200), 
        .C1(n3956), .Y(n1749) );
  OAI222XL U3372 ( .A0(n1087), .A1(n3188), .B0(n4059), .B1(n323), .C0(n4199), 
        .C1(n3956), .Y(n1748) );
  OAI222XL U3373 ( .A0(n1088), .A1(n3188), .B0(n4062), .B1(n3855), .C0(n4198), 
        .C1(n3956), .Y(n1747) );
  OAI222XL U3374 ( .A0(n1089), .A1(n3188), .B0(n4065), .B1(n3855), .C0(n4197), 
        .C1(n3956), .Y(n1746) );
  OAI222XL U3375 ( .A0(n1090), .A1(n3188), .B0(n4068), .B1(n3855), .C0(n4196), 
        .C1(n3956), .Y(n1745) );
  OAI222XL U3376 ( .A0(n1091), .A1(n3188), .B0(n4071), .B1(n3855), .C0(n4195), 
        .C1(n3956), .Y(n1744) );
  OAI222XL U3377 ( .A0(n1092), .A1(n3188), .B0(n4074), .B1(n3855), .C0(n4194), 
        .C1(n3956), .Y(n1743) );
  OAI222XL U3378 ( .A0(n1093), .A1(n3188), .B0(n4077), .B1(n3855), .C0(n4193), 
        .C1(n3956), .Y(n1742) );
  OAI222XL U3379 ( .A0(n1094), .A1(n3188), .B0(n4080), .B1(n3855), .C0(n4192), 
        .C1(n3956), .Y(n1741) );
  OAI222XL U3380 ( .A0(n1095), .A1(n3188), .B0(n4083), .B1(n3855), .C0(n4191), 
        .C1(n3956), .Y(n1740) );
  OAI222XL U3381 ( .A0(n1096), .A1(n3188), .B0(n4086), .B1(n3855), .C0(n4190), 
        .C1(n3956), .Y(n1739) );
  OAI222XL U3382 ( .A0(n1097), .A1(n3188), .B0(n4089), .B1(n3855), .C0(n4189), 
        .C1(n3956), .Y(n1738) );
  OAI222XL U3383 ( .A0(n1098), .A1(n3188), .B0(n4092), .B1(n3855), .C0(n4188), 
        .C1(n3956), .Y(n1737) );
  OAI222XL U3384 ( .A0(n1099), .A1(n3188), .B0(n4095), .B1(n3855), .C0(n4187), 
        .C1(n3949), .Y(n1736) );
  OAI222XL U3385 ( .A0(n1100), .A1(n3188), .B0(n4098), .B1(n3854), .C0(n4186), 
        .C1(n3956), .Y(n1735) );
  OAI222XL U3386 ( .A0(n1101), .A1(n3188), .B0(n4101), .B1(n3854), .C0(n4185), 
        .C1(n3949), .Y(n1734) );
  OAI222XL U3387 ( .A0(n1102), .A1(n3188), .B0(n4104), .B1(n3854), .C0(n4184), 
        .C1(n3956), .Y(n1733) );
  OAI222XL U3388 ( .A0(n1103), .A1(n3188), .B0(n4107), .B1(n3854), .C0(n4183), 
        .C1(n3955), .Y(n1732) );
  OAI222XL U3389 ( .A0(n1104), .A1(n3188), .B0(n4110), .B1(n3854), .C0(n4182), 
        .C1(n3949), .Y(n1731) );
  OAI222XL U3390 ( .A0(n1105), .A1(n3188), .B0(n4029), .B1(n3854), .C0(n4181), 
        .C1(n3951), .Y(n1730) );
  OAI222XL U3391 ( .A0(n1106), .A1(n3188), .B0(n4031), .B1(n3854), .C0(n4180), 
        .C1(n3949), .Y(n1729) );
  OAI222XL U3392 ( .A0(n1107), .A1(n3188), .B0(n4033), .B1(n3854), .C0(n4179), 
        .C1(n3955), .Y(n1728) );
  OAI222XL U3393 ( .A0(n1108), .A1(n3188), .B0(n4035), .B1(n3854), .C0(n4178), 
        .C1(n3949), .Y(n1727) );
  OAI222XL U3394 ( .A0(n1109), .A1(n3188), .B0(n4037), .B1(n3854), .C0(n4177), 
        .C1(n3949), .Y(n1726) );
  OAI222XL U3395 ( .A0(n1110), .A1(n3188), .B0(n4039), .B1(n3854), .C0(n4176), 
        .C1(n3949), .Y(n1725) );
  OAI222XL U3396 ( .A0(n1111), .A1(n3188), .B0(n4041), .B1(n3854), .C0(n4175), 
        .C1(n3951), .Y(n1724) );
  OAI222XL U3397 ( .A0(n1479), .A1(n4016), .B0(n4044), .B1(n3265), .C0(n4206), 
        .C1(n3864), .Y(n2651) );
  OAI222XL U3398 ( .A0(n1480), .A1(n4016), .B0(n4047), .B1(n3265), .C0(n4205), 
        .C1(n3864), .Y(n2650) );
  OAI222XL U3399 ( .A0(n1481), .A1(n4016), .B0(n4049), .B1(n3265), .C0(n4204), 
        .C1(n3865), .Y(n2649) );
  OAI222XL U3400 ( .A0(n1482), .A1(n4016), .B0(n4051), .B1(n3265), .C0(n4203), 
        .C1(n3865), .Y(n2648) );
  OAI222XL U3401 ( .A0(n1483), .A1(n4016), .B0(n4053), .B1(n3265), .C0(n4202), 
        .C1(n3865), .Y(n2647) );
  OAI222XL U3402 ( .A0(n1484), .A1(n4016), .B0(n4055), .B1(n3265), .C0(n4201), 
        .C1(n3865), .Y(n2646) );
  OAI222XL U3403 ( .A0(n1485), .A1(n4016), .B0(n4057), .B1(n3265), .C0(n4200), 
        .C1(n3865), .Y(n2645) );
  OAI222XL U3404 ( .A0(n1486), .A1(n4016), .B0(n4059), .B1(n3265), .C0(n4199), 
        .C1(n3865), .Y(n2644) );
  OAI222XL U3405 ( .A0(n1487), .A1(n4016), .B0(n4062), .B1(n3265), .C0(n4198), 
        .C1(n3865), .Y(n2643) );
  OAI222XL U3406 ( .A0(n1488), .A1(n4016), .B0(n4065), .B1(n3265), .C0(n4197), 
        .C1(n3865), .Y(n2642) );
  OAI222XL U3407 ( .A0(n1489), .A1(n4016), .B0(n4068), .B1(n3265), .C0(n4196), 
        .C1(n3865), .Y(n2641) );
  OAI222XL U3408 ( .A0(n1490), .A1(n4016), .B0(n4071), .B1(n3265), .C0(n4195), 
        .C1(n3865), .Y(n2640) );
  OAI222XL U3409 ( .A0(n1491), .A1(n4016), .B0(n4074), .B1(n3265), .C0(n4194), 
        .C1(n3865), .Y(n2639) );
  OAI222XL U3410 ( .A0(n1492), .A1(n4016), .B0(n4077), .B1(n3265), .C0(n4193), 
        .C1(n3865), .Y(n2638) );
  OAI222XL U3411 ( .A0(n1493), .A1(n4016), .B0(n4080), .B1(n3265), .C0(n4192), 
        .C1(n3865), .Y(n2637) );
  OAI222XL U3412 ( .A0(n1494), .A1(n4016), .B0(n4083), .B1(n3265), .C0(n4191), 
        .C1(n3865), .Y(n2636) );
  OAI222XL U3413 ( .A0(n1495), .A1(n4016), .B0(n4086), .B1(n3265), .C0(n4190), 
        .C1(n3865), .Y(n2635) );
  OAI222XL U3414 ( .A0(n1496), .A1(n4016), .B0(n4089), .B1(n3265), .C0(n4189), 
        .C1(n3865), .Y(n2634) );
  OAI222XL U3415 ( .A0(n1497), .A1(n4016), .B0(n4092), .B1(n3265), .C0(n4188), 
        .C1(n3859), .Y(n2633) );
  OAI222XL U3416 ( .A0(n1498), .A1(n4016), .B0(n4095), .B1(n3265), .C0(n4187), 
        .C1(n3859), .Y(n2632) );
  OAI222XL U3417 ( .A0(n1499), .A1(n4016), .B0(n4098), .B1(n3265), .C0(n4186), 
        .C1(n3859), .Y(n2631) );
  OAI222XL U3418 ( .A0(n1500), .A1(n4016), .B0(n4101), .B1(n3265), .C0(n4185), 
        .C1(n3858), .Y(n2630) );
  OAI222XL U3419 ( .A0(n1501), .A1(n4016), .B0(n4104), .B1(n3265), .C0(n4184), 
        .C1(n3859), .Y(n2629) );
  OAI222XL U3420 ( .A0(n1502), .A1(n4016), .B0(n4107), .B1(n3265), .C0(n4183), 
        .C1(n3858), .Y(n2628) );
  OAI222XL U3421 ( .A0(n1503), .A1(n4016), .B0(n4110), .B1(n3265), .C0(n4182), 
        .C1(n3859), .Y(n2627) );
  OAI222XL U3422 ( .A0(n1504), .A1(n4016), .B0(n3214), .B1(n3265), .C0(n4181), 
        .C1(n3858), .Y(n2626) );
  OAI222XL U3423 ( .A0(n1505), .A1(n4016), .B0(n3215), .B1(n3265), .C0(n4180), 
        .C1(n3859), .Y(n2625) );
  OAI222XL U3424 ( .A0(n1506), .A1(n4016), .B0(n3216), .B1(n3265), .C0(n4179), 
        .C1(n3862), .Y(n2624) );
  OAI222XL U3425 ( .A0(n1507), .A1(n4016), .B0(n3205), .B1(n3265), .C0(n4178), 
        .C1(n3858), .Y(n2623) );
  OAI222XL U3426 ( .A0(n1508), .A1(n4016), .B0(n3206), .B1(n3265), .C0(n4177), 
        .C1(n3859), .Y(n2622) );
  OAI222XL U3427 ( .A0(n1509), .A1(n4016), .B0(n3207), .B1(n3265), .C0(n4176), 
        .C1(n3861), .Y(n2621) );
  OAI222XL U3428 ( .A0(n1510), .A1(n4016), .B0(n3208), .B1(n3265), .C0(n4175), 
        .C1(n3864), .Y(n2620) );
  OAI222XL U3429 ( .A0(n1607), .A1(n4027), .B0(n4044), .B1(n3184), .C0(n3878), 
        .C1(n4206), .Y(n2523) );
  OAI222XL U3430 ( .A0(n1608), .A1(n4027), .B0(n4047), .B1(n3184), .C0(n3878), 
        .C1(n4205), .Y(n2522) );
  OAI222XL U3431 ( .A0(n1609), .A1(n4027), .B0(n4049), .B1(n3184), .C0(n3878), 
        .C1(n4204), .Y(n2521) );
  OAI222XL U3432 ( .A0(n1610), .A1(n4027), .B0(n4051), .B1(n3184), .C0(n3878), 
        .C1(n4203), .Y(n2520) );
  OAI222XL U3433 ( .A0(n1611), .A1(n4027), .B0(n4053), .B1(n3184), .C0(n3879), 
        .C1(n4202), .Y(n2519) );
  OAI222XL U3434 ( .A0(n1612), .A1(n4027), .B0(n4055), .B1(n3184), .C0(n3879), 
        .C1(n4201), .Y(n2518) );
  OAI222XL U3435 ( .A0(n1613), .A1(n4027), .B0(n4057), .B1(n3184), .C0(n3879), 
        .C1(n4200), .Y(n2517) );
  OAI222XL U3436 ( .A0(n1614), .A1(n4027), .B0(n4059), .B1(n3184), .C0(n3879), 
        .C1(n4199), .Y(n2516) );
  OAI222XL U3437 ( .A0(n1615), .A1(n4027), .B0(n4062), .B1(n3184), .C0(n3879), 
        .C1(n4198), .Y(n2515) );
  OAI222XL U3438 ( .A0(n1616), .A1(n4027), .B0(n4065), .B1(n3184), .C0(n3879), 
        .C1(n4197), .Y(n2514) );
  OAI222XL U3439 ( .A0(n1617), .A1(n4027), .B0(n4068), .B1(n3184), .C0(n3879), 
        .C1(n4196), .Y(n2513) );
  OAI222XL U3440 ( .A0(n1618), .A1(n4027), .B0(n4071), .B1(n3184), .C0(n3879), 
        .C1(n4195), .Y(n2512) );
  OAI222XL U3441 ( .A0(n1619), .A1(n4027), .B0(n4074), .B1(n3184), .C0(n3879), 
        .C1(n4194), .Y(n2511) );
  OAI222XL U3442 ( .A0(n1620), .A1(n4027), .B0(n4077), .B1(n3184), .C0(n3879), 
        .C1(n4193), .Y(n2510) );
  OAI222XL U3443 ( .A0(n1621), .A1(n4027), .B0(n4080), .B1(n3184), .C0(n3879), 
        .C1(n4192), .Y(n2509) );
  OAI222XL U3444 ( .A0(n1622), .A1(n4027), .B0(n4083), .B1(n3184), .C0(n3879), 
        .C1(n4191), .Y(n2508) );
  OAI222XL U3445 ( .A0(n1623), .A1(n4027), .B0(n4086), .B1(n3184), .C0(n3879), 
        .C1(n4190), .Y(n2507) );
  OAI222XL U3446 ( .A0(n1624), .A1(n4027), .B0(n4089), .B1(n3184), .C0(n3879), 
        .C1(n4189), .Y(n2506) );
  OAI222XL U3447 ( .A0(n1625), .A1(n4027), .B0(n4092), .B1(n3184), .C0(n3879), 
        .C1(n4188), .Y(n2505) );
  OAI222XL U3448 ( .A0(n1626), .A1(n4027), .B0(n4095), .B1(n3184), .C0(n3879), 
        .C1(n4187), .Y(n2504) );
  OAI222XL U3449 ( .A0(n1627), .A1(n4027), .B0(n4098), .B1(n3184), .C0(n3871), 
        .C1(n4186), .Y(n2503) );
  OAI222XL U3450 ( .A0(n1628), .A1(n4027), .B0(n4101), .B1(n3184), .C0(n3879), 
        .C1(n4185), .Y(n2502) );
  OAI222XL U3451 ( .A0(n1629), .A1(n4027), .B0(n4104), .B1(n3184), .C0(n3871), 
        .C1(n4184), .Y(n2501) );
  OAI222XL U3452 ( .A0(n1630), .A1(n4027), .B0(n4107), .B1(n3184), .C0(n3879), 
        .C1(n4183), .Y(n2500) );
  OAI222XL U3453 ( .A0(n1631), .A1(n4027), .B0(n4110), .B1(n3184), .C0(n3879), 
        .C1(n4182), .Y(n2499) );
  OAI222XL U3454 ( .A0(n1632), .A1(n4027), .B0(n4028), .B1(n3184), .C0(n3871), 
        .C1(n4181), .Y(n2498) );
  OAI222XL U3455 ( .A0(n1633), .A1(n4027), .B0(n4030), .B1(n3184), .C0(n3871), 
        .C1(n4180), .Y(n2497) );
  OAI222XL U3456 ( .A0(n1634), .A1(n4027), .B0(n4032), .B1(n3184), .C0(n3879), 
        .C1(n4179), .Y(n2496) );
  OAI222XL U3457 ( .A0(n1635), .A1(n4027), .B0(n4034), .B1(n3184), .C0(n3874), 
        .C1(n4178), .Y(n2495) );
  OAI222XL U3458 ( .A0(n1636), .A1(n4027), .B0(n4036), .B1(n3184), .C0(n3871), 
        .C1(n4177), .Y(n2494) );
  OAI222XL U3459 ( .A0(n1637), .A1(n4027), .B0(n4038), .B1(n3184), .C0(n3873), 
        .C1(n4176), .Y(n2493) );
  OAI222XL U3460 ( .A0(n1638), .A1(n4027), .B0(n4040), .B1(n3184), .C0(n3871), 
        .C1(n4175), .Y(n2492) );
  OAI222XL U3461 ( .A0(n472), .A1(n3198), .B0(n4043), .B1(n3817), .C0(n4302), 
        .C1(n3898), .Y(n2363) );
  OAI222XL U3462 ( .A0(n473), .A1(n3198), .B0(n4046), .B1(n3816), .C0(n4301), 
        .C1(n3899), .Y(n2362) );
  OAI222XL U3463 ( .A0(n474), .A1(n3198), .B0(n4049), .B1(n361), .C0(n4300), 
        .C1(n3898), .Y(n2361) );
  OAI222XL U3464 ( .A0(n475), .A1(n3198), .B0(n4051), .B1(n361), .C0(n4299), 
        .C1(n3899), .Y(n2360) );
  OAI222XL U3465 ( .A0(n476), .A1(n3198), .B0(n4053), .B1(n361), .C0(n4298), 
        .C1(n3899), .Y(n2359) );
  OAI222XL U3466 ( .A0(n477), .A1(n3198), .B0(n4055), .B1(n361), .C0(n4297), 
        .C1(n3898), .Y(n2358) );
  OAI222XL U3467 ( .A0(n478), .A1(n3198), .B0(n4057), .B1(n361), .C0(n4296), 
        .C1(n3898), .Y(n2357) );
  OAI222XL U3468 ( .A0(n479), .A1(n3198), .B0(n4059), .B1(n361), .C0(n4295), 
        .C1(n3899), .Y(n2356) );
  OAI222XL U3469 ( .A0(n480), .A1(n3198), .B0(n4061), .B1(n3817), .C0(n4294), 
        .C1(n3899), .Y(n2355) );
  OAI222XL U3470 ( .A0(n481), .A1(n3198), .B0(n4064), .B1(n3817), .C0(n4293), 
        .C1(n3899), .Y(n2354) );
  OAI222XL U3471 ( .A0(n482), .A1(n3198), .B0(n4067), .B1(n3817), .C0(n4292), 
        .C1(n3899), .Y(n2353) );
  OAI222XL U3472 ( .A0(n483), .A1(n3198), .B0(n4070), .B1(n3817), .C0(n4291), 
        .C1(n3904), .Y(n2352) );
  OAI222XL U3473 ( .A0(n484), .A1(n3198), .B0(n4073), .B1(n3817), .C0(n4290), 
        .C1(n3899), .Y(n2351) );
  OAI222XL U3474 ( .A0(n485), .A1(n3198), .B0(n4076), .B1(n3817), .C0(n4289), 
        .C1(n3899), .Y(n2350) );
  OAI222XL U3475 ( .A0(n486), .A1(n3198), .B0(n4079), .B1(n3817), .C0(n4288), 
        .C1(n3899), .Y(n2349) );
  OAI222XL U3476 ( .A0(n487), .A1(n3198), .B0(n4082), .B1(n3817), .C0(n4287), 
        .C1(n3899), .Y(n2348) );
  OAI222XL U3477 ( .A0(n488), .A1(n3198), .B0(n4085), .B1(n3817), .C0(n4286), 
        .C1(n3899), .Y(n2347) );
  OAI222XL U3478 ( .A0(n489), .A1(n3198), .B0(n4088), .B1(n3817), .C0(n4285), 
        .C1(n3899), .Y(n2346) );
  OAI222XL U3479 ( .A0(n490), .A1(n3198), .B0(n4091), .B1(n3817), .C0(n4284), 
        .C1(n3899), .Y(n2345) );
  OAI222XL U3480 ( .A0(n491), .A1(n3198), .B0(n4094), .B1(n3817), .C0(n4283), 
        .C1(n3901), .Y(n2344) );
  OAI222XL U3481 ( .A0(n492), .A1(n3198), .B0(n4097), .B1(n3816), .C0(n4282), 
        .C1(n3899), .Y(n2343) );
  OAI222XL U3482 ( .A0(n493), .A1(n3198), .B0(n4100), .B1(n3816), .C0(n4281), 
        .C1(n3899), .Y(n2342) );
  OAI222XL U3483 ( .A0(n494), .A1(n3198), .B0(n4103), .B1(n3816), .C0(n4280), 
        .C1(n3902), .Y(n2341) );
  OAI222XL U3484 ( .A0(n495), .A1(n3198), .B0(n4106), .B1(n3816), .C0(n4279), 
        .C1(n3899), .Y(n2340) );
  OAI222XL U3485 ( .A0(n496), .A1(n3198), .B0(n3209), .B1(n3816), .C0(n4278), 
        .C1(n3903), .Y(n2339) );
  OAI222XL U3486 ( .A0(n497), .A1(n3198), .B0(n4028), .B1(n3816), .C0(n4277), 
        .C1(n3903), .Y(n2338) );
  OAI222XL U3487 ( .A0(n498), .A1(n3198), .B0(n4030), .B1(n3816), .C0(n4276), 
        .C1(n3899), .Y(n2337) );
  OAI222XL U3488 ( .A0(n499), .A1(n3198), .B0(n4032), .B1(n3816), .C0(n4275), 
        .C1(n3900), .Y(n2336) );
  OAI222XL U3489 ( .A0(n500), .A1(n3198), .B0(n4034), .B1(n3816), .C0(n4274), 
        .C1(n3897), .Y(n2335) );
  OAI222XL U3490 ( .A0(n501), .A1(n3198), .B0(n4036), .B1(n3816), .C0(n4273), 
        .C1(n3903), .Y(n2334) );
  OAI222XL U3491 ( .A0(n502), .A1(n3198), .B0(n4038), .B1(n3816), .C0(n4272), 
        .C1(n3897), .Y(n2333) );
  OAI222XL U3492 ( .A0(n503), .A1(n3198), .B0(n4040), .B1(n3816), .C0(n4271), 
        .C1(n3904), .Y(n2332) );
  OAI222XL U3493 ( .A0(n600), .A1(n3197), .B0(n4045), .B1(n3825), .C0(n4302), 
        .C1(n3911), .Y(n2235) );
  OAI222XL U3494 ( .A0(n601), .A1(n3197), .B0(n4048), .B1(n3824), .C0(n4301), 
        .C1(n3912), .Y(n2234) );
  OAI222XL U3495 ( .A0(n602), .A1(n3197), .B0(n4050), .B1(n353), .C0(n4300), 
        .C1(n3911), .Y(n2233) );
  OAI222XL U3496 ( .A0(n603), .A1(n3197), .B0(n4052), .B1(n353), .C0(n4299), 
        .C1(n3912), .Y(n2232) );
  OAI222XL U3497 ( .A0(n604), .A1(n3197), .B0(n4054), .B1(n353), .C0(n4298), 
        .C1(n3912), .Y(n2231) );
  OAI222XL U3498 ( .A0(n605), .A1(n3197), .B0(n4056), .B1(n353), .C0(n4297), 
        .C1(n3911), .Y(n2230) );
  OAI222XL U3499 ( .A0(n606), .A1(n3197), .B0(n4058), .B1(n353), .C0(n4296), 
        .C1(n3911), .Y(n2229) );
  OAI222XL U3500 ( .A0(n607), .A1(n3197), .B0(n4060), .B1(n353), .C0(n4295), 
        .C1(n3912), .Y(n2228) );
  OAI222XL U3501 ( .A0(n608), .A1(n3197), .B0(n4063), .B1(n3825), .C0(n4294), 
        .C1(n3912), .Y(n2227) );
  OAI222XL U3502 ( .A0(n609), .A1(n3197), .B0(n4066), .B1(n3825), .C0(n4293), 
        .C1(n3912), .Y(n2226) );
  OAI222XL U3503 ( .A0(n610), .A1(n3197), .B0(n4069), .B1(n3825), .C0(n4292), 
        .C1(n3912), .Y(n2225) );
  OAI222XL U3504 ( .A0(n611), .A1(n3197), .B0(n4072), .B1(n3825), .C0(n4291), 
        .C1(n3912), .Y(n2224) );
  OAI222XL U3505 ( .A0(n612), .A1(n3197), .B0(n4075), .B1(n3825), .C0(n4290), 
        .C1(n3912), .Y(n2223) );
  OAI222XL U3506 ( .A0(n613), .A1(n3197), .B0(n4078), .B1(n3825), .C0(n4289), 
        .C1(n3916), .Y(n2222) );
  OAI222XL U3507 ( .A0(n614), .A1(n3197), .B0(n4081), .B1(n3825), .C0(n4288), 
        .C1(n3912), .Y(n2221) );
  OAI222XL U3508 ( .A0(n615), .A1(n3197), .B0(n4084), .B1(n3825), .C0(n4287), 
        .C1(n3912), .Y(n2220) );
  OAI222XL U3509 ( .A0(n616), .A1(n3197), .B0(n4087), .B1(n3825), .C0(n4286), 
        .C1(n3913), .Y(n2219) );
  OAI222XL U3510 ( .A0(n617), .A1(n3197), .B0(n4090), .B1(n3825), .C0(n4285), 
        .C1(n3912), .Y(n2218) );
  OAI222XL U3511 ( .A0(n618), .A1(n3197), .B0(n4093), .B1(n3825), .C0(n4284), 
        .C1(n3912), .Y(n2217) );
  OAI222XL U3512 ( .A0(n619), .A1(n3197), .B0(n4096), .B1(n3825), .C0(n4283), 
        .C1(n3914), .Y(n2216) );
  OAI222XL U3513 ( .A0(n620), .A1(n3197), .B0(n4099), .B1(n3824), .C0(n4282), 
        .C1(n3912), .Y(n2215) );
  OAI222XL U3514 ( .A0(n621), .A1(n3197), .B0(n4102), .B1(n3824), .C0(n4281), 
        .C1(n3912), .Y(n2214) );
  OAI222XL U3515 ( .A0(n622), .A1(n3197), .B0(n4105), .B1(n3824), .C0(n4280), 
        .C1(n3915), .Y(n2213) );
  OAI222XL U3516 ( .A0(n623), .A1(n3197), .B0(n4108), .B1(n3824), .C0(n4279), 
        .C1(n3912), .Y(n2212) );
  OAI222XL U3517 ( .A0(n624), .A1(n3197), .B0(n3209), .B1(n3824), .C0(n4278), 
        .C1(n3917), .Y(n2211) );
  OAI222XL U3518 ( .A0(n625), .A1(n3197), .B0(n4028), .B1(n3824), .C0(n4277), 
        .C1(n3914), .Y(n2210) );
  OAI222XL U3519 ( .A0(n626), .A1(n3197), .B0(n4030), .B1(n3824), .C0(n4276), 
        .C1(n3916), .Y(n2209) );
  OAI222XL U3520 ( .A0(n627), .A1(n3197), .B0(n4032), .B1(n3824), .C0(n4275), 
        .C1(n3915), .Y(n2208) );
  OAI222XL U3521 ( .A0(n628), .A1(n3197), .B0(n4034), .B1(n3824), .C0(n4274), 
        .C1(n3917), .Y(n2207) );
  OAI222XL U3522 ( .A0(n629), .A1(n3197), .B0(n4036), .B1(n3824), .C0(n4273), 
        .C1(n3913), .Y(n2206) );
  OAI222XL U3523 ( .A0(n630), .A1(n3197), .B0(n4038), .B1(n3824), .C0(n4272), 
        .C1(n3912), .Y(n2205) );
  OAI222XL U3524 ( .A0(n631), .A1(n3197), .B0(n4040), .B1(n3824), .C0(n4271), 
        .C1(n3916), .Y(n2204) );
  OAI222XL U3525 ( .A0(n728), .A1(n3196), .B0(n4045), .B1(n3833), .C0(n4302), 
        .C1(n3924), .Y(n2107) );
  OAI222XL U3526 ( .A0(n729), .A1(n3196), .B0(n4048), .B1(n3832), .C0(n4301), 
        .C1(n3925), .Y(n2106) );
  OAI222XL U3527 ( .A0(n730), .A1(n3196), .B0(n4050), .B1(n345), .C0(n4300), 
        .C1(n3924), .Y(n2105) );
  OAI222XL U3528 ( .A0(n731), .A1(n3196), .B0(n4052), .B1(n345), .C0(n4299), 
        .C1(n3925), .Y(n2104) );
  OAI222XL U3529 ( .A0(n732), .A1(n3196), .B0(n4054), .B1(n345), .C0(n4298), 
        .C1(n3925), .Y(n2103) );
  OAI222XL U3530 ( .A0(n733), .A1(n3196), .B0(n4056), .B1(n345), .C0(n4297), 
        .C1(n3924), .Y(n2102) );
  OAI222XL U3531 ( .A0(n734), .A1(n3196), .B0(n4058), .B1(n345), .C0(n4296), 
        .C1(n3924), .Y(n2101) );
  OAI222XL U3532 ( .A0(n735), .A1(n3196), .B0(n4060), .B1(n345), .C0(n4295), 
        .C1(n3925), .Y(n2100) );
  OAI222XL U3533 ( .A0(n736), .A1(n3196), .B0(n4063), .B1(n3833), .C0(n4294), 
        .C1(n3925), .Y(n2099) );
  OAI222XL U3534 ( .A0(n737), .A1(n3196), .B0(n4066), .B1(n3833), .C0(n4293), 
        .C1(n3925), .Y(n2098) );
  OAI222XL U3535 ( .A0(n738), .A1(n3196), .B0(n4069), .B1(n3833), .C0(n4292), 
        .C1(n3925), .Y(n2097) );
  OAI222XL U3536 ( .A0(n739), .A1(n3196), .B0(n4072), .B1(n3833), .C0(n4291), 
        .C1(n3925), .Y(n2096) );
  OAI222XL U3537 ( .A0(n740), .A1(n3196), .B0(n4075), .B1(n3833), .C0(n4290), 
        .C1(n3925), .Y(n2095) );
  OAI222XL U3538 ( .A0(n741), .A1(n3196), .B0(n4078), .B1(n3833), .C0(n4289), 
        .C1(n3929), .Y(n2094) );
  OAI222XL U3539 ( .A0(n742), .A1(n3196), .B0(n4081), .B1(n3833), .C0(n4288), 
        .C1(n3925), .Y(n2093) );
  OAI222XL U3540 ( .A0(n743), .A1(n3196), .B0(n4084), .B1(n3833), .C0(n4287), 
        .C1(n3925), .Y(n2092) );
  OAI222XL U3541 ( .A0(n744), .A1(n3196), .B0(n4087), .B1(n3833), .C0(n4286), 
        .C1(n3926), .Y(n2091) );
  OAI222XL U3542 ( .A0(n745), .A1(n3196), .B0(n4090), .B1(n3833), .C0(n4285), 
        .C1(n3925), .Y(n2090) );
  OAI222XL U3543 ( .A0(n746), .A1(n3196), .B0(n4093), .B1(n3833), .C0(n4284), 
        .C1(n3925), .Y(n2089) );
  OAI222XL U3544 ( .A0(n747), .A1(n3196), .B0(n4096), .B1(n3833), .C0(n4283), 
        .C1(n3927), .Y(n2088) );
  OAI222XL U3545 ( .A0(n748), .A1(n3196), .B0(n4099), .B1(n3832), .C0(n4282), 
        .C1(n3925), .Y(n2087) );
  OAI222XL U3546 ( .A0(n749), .A1(n3196), .B0(n4102), .B1(n3832), .C0(n4281), 
        .C1(n3925), .Y(n2086) );
  OAI222XL U3547 ( .A0(n750), .A1(n3196), .B0(n4105), .B1(n3832), .C0(n4280), 
        .C1(n3928), .Y(n2085) );
  OAI222XL U3548 ( .A0(n751), .A1(n3196), .B0(n4108), .B1(n3832), .C0(n4279), 
        .C1(n3925), .Y(n2084) );
  OAI222XL U3549 ( .A0(n752), .A1(n3196), .B0(n4111), .B1(n3832), .C0(n4278), 
        .C1(n3930), .Y(n2083) );
  OAI222XL U3550 ( .A0(n753), .A1(n3196), .B0(n4028), .B1(n3832), .C0(n4277), 
        .C1(n3927), .Y(n2082) );
  OAI222XL U3551 ( .A0(n754), .A1(n3196), .B0(n4030), .B1(n3832), .C0(n4276), 
        .C1(n3929), .Y(n2081) );
  OAI222XL U3552 ( .A0(n755), .A1(n3196), .B0(n4032), .B1(n3832), .C0(n4275), 
        .C1(n3928), .Y(n2080) );
  OAI222XL U3553 ( .A0(n756), .A1(n3196), .B0(n4034), .B1(n3832), .C0(n4274), 
        .C1(n3930), .Y(n2079) );
  OAI222XL U3554 ( .A0(n757), .A1(n3196), .B0(n4036), .B1(n3832), .C0(n4273), 
        .C1(n3926), .Y(n2078) );
  OAI222XL U3555 ( .A0(n758), .A1(n3196), .B0(n4038), .B1(n3832), .C0(n4272), 
        .C1(n3925), .Y(n2077) );
  OAI222XL U3556 ( .A0(n759), .A1(n3196), .B0(n4040), .B1(n3832), .C0(n4271), 
        .C1(n3929), .Y(n2076) );
  OAI222XL U3557 ( .A0(n856), .A1(n3199), .B0(n4045), .B1(n3841), .C0(n4302), 
        .C1(n3937), .Y(n1979) );
  OAI222XL U3558 ( .A0(n857), .A1(n3199), .B0(n4048), .B1(n3840), .C0(n4301), 
        .C1(n3938), .Y(n1978) );
  OAI222XL U3559 ( .A0(n858), .A1(n3199), .B0(n4050), .B1(n337), .C0(n4300), 
        .C1(n3937), .Y(n1977) );
  OAI222XL U3560 ( .A0(n859), .A1(n3199), .B0(n4052), .B1(n337), .C0(n4299), 
        .C1(n3938), .Y(n1976) );
  OAI222XL U3561 ( .A0(n860), .A1(n3199), .B0(n4054), .B1(n337), .C0(n4298), 
        .C1(n3938), .Y(n1975) );
  OAI222XL U3562 ( .A0(n861), .A1(n3199), .B0(n4056), .B1(n337), .C0(n4297), 
        .C1(n3937), .Y(n1974) );
  OAI222XL U3563 ( .A0(n862), .A1(n3199), .B0(n4058), .B1(n337), .C0(n4296), 
        .C1(n3937), .Y(n1973) );
  OAI222XL U3564 ( .A0(n863), .A1(n3199), .B0(n4060), .B1(n337), .C0(n4295), 
        .C1(n3938), .Y(n1972) );
  OAI222XL U3565 ( .A0(n864), .A1(n3199), .B0(n4063), .B1(n3841), .C0(n4294), 
        .C1(n3938), .Y(n1971) );
  OAI222XL U3566 ( .A0(n865), .A1(n3199), .B0(n4066), .B1(n3841), .C0(n4293), 
        .C1(n3938), .Y(n1970) );
  OAI222XL U3567 ( .A0(n866), .A1(n3199), .B0(n4069), .B1(n3841), .C0(n4292), 
        .C1(n3938), .Y(n1969) );
  OAI222XL U3568 ( .A0(n867), .A1(n3199), .B0(n4072), .B1(n3841), .C0(n4291), 
        .C1(n3938), .Y(n1968) );
  OAI222XL U3569 ( .A0(n868), .A1(n3199), .B0(n4075), .B1(n3841), .C0(n4290), 
        .C1(n3938), .Y(n1967) );
  OAI222XL U3570 ( .A0(n869), .A1(n3199), .B0(n4078), .B1(n3841), .C0(n4289), 
        .C1(n3942), .Y(n1966) );
  OAI222XL U3571 ( .A0(n870), .A1(n3199), .B0(n4081), .B1(n3841), .C0(n4288), 
        .C1(n3938), .Y(n1965) );
  OAI222XL U3572 ( .A0(n871), .A1(n3199), .B0(n4084), .B1(n3841), .C0(n4287), 
        .C1(n3938), .Y(n1964) );
  OAI222XL U3573 ( .A0(n872), .A1(n3199), .B0(n4087), .B1(n3841), .C0(n4286), 
        .C1(n3939), .Y(n1963) );
  OAI222XL U3574 ( .A0(n873), .A1(n3199), .B0(n4090), .B1(n3841), .C0(n4285), 
        .C1(n3938), .Y(n1962) );
  OAI222XL U3575 ( .A0(n874), .A1(n3199), .B0(n4093), .B1(n3841), .C0(n4284), 
        .C1(n3938), .Y(n1961) );
  OAI222XL U3576 ( .A0(n875), .A1(n3199), .B0(n4096), .B1(n3841), .C0(n4283), 
        .C1(n3940), .Y(n1960) );
  OAI222XL U3577 ( .A0(n876), .A1(n3199), .B0(n4099), .B1(n3840), .C0(n4282), 
        .C1(n3938), .Y(n1959) );
  OAI222XL U3578 ( .A0(n877), .A1(n3199), .B0(n4102), .B1(n3840), .C0(n4281), 
        .C1(n3938), .Y(n1958) );
  OAI222XL U3579 ( .A0(n878), .A1(n3199), .B0(n4105), .B1(n3840), .C0(n4280), 
        .C1(n3941), .Y(n1957) );
  OAI222XL U3580 ( .A0(n879), .A1(n3199), .B0(n4108), .B1(n3840), .C0(n4279), 
        .C1(n3938), .Y(n1956) );
  OAI222XL U3581 ( .A0(n880), .A1(n3199), .B0(n4111), .B1(n3840), .C0(n4278), 
        .C1(n3943), .Y(n1955) );
  OAI222XL U3582 ( .A0(n881), .A1(n3199), .B0(n4029), .B1(n3840), .C0(n4277), 
        .C1(n3942), .Y(n1954) );
  OAI222XL U3583 ( .A0(n882), .A1(n3199), .B0(n4031), .B1(n3840), .C0(n4276), 
        .C1(n3939), .Y(n1953) );
  OAI222XL U3584 ( .A0(n883), .A1(n3199), .B0(n4033), .B1(n3840), .C0(n4275), 
        .C1(n3940), .Y(n1952) );
  OAI222XL U3585 ( .A0(n884), .A1(n3199), .B0(n4035), .B1(n3840), .C0(n4274), 
        .C1(n3936), .Y(n1951) );
  OAI222XL U3586 ( .A0(n885), .A1(n3199), .B0(n4037), .B1(n3840), .C0(n4273), 
        .C1(n3941), .Y(n1950) );
  OAI222XL U3587 ( .A0(n886), .A1(n3199), .B0(n4039), .B1(n3840), .C0(n4272), 
        .C1(n3943), .Y(n1949) );
  OAI222XL U3588 ( .A0(n887), .A1(n3199), .B0(n4041), .B1(n3840), .C0(n4271), 
        .C1(n3938), .Y(n1948) );
  OAI222XL U3589 ( .A0(n984), .A1(n3200), .B0(n4045), .B1(n3849), .C0(n4302), 
        .C1(n3950), .Y(n1851) );
  OAI222XL U3590 ( .A0(n985), .A1(n3200), .B0(n4048), .B1(n3848), .C0(n4301), 
        .C1(n3951), .Y(n1850) );
  OAI222XL U3591 ( .A0(n986), .A1(n3200), .B0(n4050), .B1(n329), .C0(n4300), 
        .C1(n3950), .Y(n1849) );
  OAI222XL U3592 ( .A0(n987), .A1(n3200), .B0(n4052), .B1(n329), .C0(n4299), 
        .C1(n3951), .Y(n1848) );
  OAI222XL U3593 ( .A0(n988), .A1(n3200), .B0(n4054), .B1(n329), .C0(n4298), 
        .C1(n3951), .Y(n1847) );
  OAI222XL U3594 ( .A0(n989), .A1(n3200), .B0(n4056), .B1(n329), .C0(n4297), 
        .C1(n3950), .Y(n1846) );
  OAI222XL U3595 ( .A0(n990), .A1(n3200), .B0(n4058), .B1(n329), .C0(n4296), 
        .C1(n3950), .Y(n1845) );
  OAI222XL U3596 ( .A0(n991), .A1(n3200), .B0(n4060), .B1(n329), .C0(n4295), 
        .C1(n3951), .Y(n1844) );
  OAI222XL U3597 ( .A0(n992), .A1(n3200), .B0(n4063), .B1(n3849), .C0(n4294), 
        .C1(n3951), .Y(n1843) );
  OAI222XL U3598 ( .A0(n993), .A1(n3200), .B0(n4066), .B1(n3849), .C0(n4293), 
        .C1(n3951), .Y(n1842) );
  OAI222XL U3599 ( .A0(n994), .A1(n3200), .B0(n4069), .B1(n3849), .C0(n4292), 
        .C1(n3951), .Y(n1841) );
  OAI222XL U3600 ( .A0(n995), .A1(n3200), .B0(n4072), .B1(n3849), .C0(n4291), 
        .C1(n3951), .Y(n1840) );
  OAI222XL U3601 ( .A0(n996), .A1(n3200), .B0(n4075), .B1(n3849), .C0(n4290), 
        .C1(n3951), .Y(n1839) );
  OAI222XL U3602 ( .A0(n997), .A1(n3200), .B0(n4078), .B1(n3849), .C0(n4289), 
        .C1(n3955), .Y(n1838) );
  OAI222XL U3603 ( .A0(n998), .A1(n3200), .B0(n4081), .B1(n3849), .C0(n4288), 
        .C1(n3951), .Y(n1837) );
  OAI222XL U3604 ( .A0(n999), .A1(n3200), .B0(n4084), .B1(n3849), .C0(n4287), 
        .C1(n3951), .Y(n1836) );
  OAI222XL U3605 ( .A0(n1000), .A1(n3200), .B0(n4087), .B1(n3849), .C0(n4286), 
        .C1(n3952), .Y(n1835) );
  OAI222XL U3606 ( .A0(n1001), .A1(n3200), .B0(n4090), .B1(n3849), .C0(n4285), 
        .C1(n3951), .Y(n1834) );
  OAI222XL U3607 ( .A0(n1002), .A1(n3200), .B0(n4093), .B1(n3849), .C0(n4284), 
        .C1(n3951), .Y(n1833) );
  OAI222XL U3608 ( .A0(n1003), .A1(n3200), .B0(n4096), .B1(n3849), .C0(n4283), 
        .C1(n3953), .Y(n1832) );
  OAI222XL U3609 ( .A0(n1004), .A1(n3200), .B0(n4099), .B1(n3848), .C0(n4282), 
        .C1(n3951), .Y(n1831) );
  OAI222XL U3610 ( .A0(n1005), .A1(n3200), .B0(n4102), .B1(n3848), .C0(n4281), 
        .C1(n3951), .Y(n1830) );
  OAI222XL U3611 ( .A0(n1006), .A1(n3200), .B0(n4105), .B1(n3848), .C0(n4280), 
        .C1(n3954), .Y(n1829) );
  OAI222XL U3612 ( .A0(n1007), .A1(n3200), .B0(n4108), .B1(n3848), .C0(n4279), 
        .C1(n3951), .Y(n1828) );
  OAI222XL U3613 ( .A0(n1008), .A1(n3200), .B0(n4111), .B1(n3848), .C0(n4278), 
        .C1(n3956), .Y(n1827) );
  OAI222XL U3614 ( .A0(n1009), .A1(n3200), .B0(n4029), .B1(n3848), .C0(n4277), 
        .C1(n3951), .Y(n1826) );
  OAI222XL U3615 ( .A0(n1010), .A1(n3200), .B0(n4031), .B1(n3848), .C0(n4276), 
        .C1(n3955), .Y(n1825) );
  OAI222XL U3616 ( .A0(n1011), .A1(n3200), .B0(n4033), .B1(n3848), .C0(n4275), 
        .C1(n3955), .Y(n1824) );
  OAI222XL U3617 ( .A0(n1012), .A1(n3200), .B0(n4035), .B1(n3848), .C0(n4274), 
        .C1(n3949), .Y(n1823) );
  OAI222XL U3618 ( .A0(n1013), .A1(n3200), .B0(n4037), .B1(n3848), .C0(n4273), 
        .C1(n3952), .Y(n1822) );
  OAI222XL U3619 ( .A0(n1014), .A1(n3200), .B0(n4039), .B1(n3848), .C0(n4272), 
        .C1(n3949), .Y(n1821) );
  OAI222XL U3620 ( .A0(n1015), .A1(n3200), .B0(n4041), .B1(n3848), .C0(n4271), 
        .C1(n3956), .Y(n1820) );
  OAI222XL U3621 ( .A0(n1383), .A1(n4009), .B0(n4044), .B1(n4006), .C0(n4302), 
        .C1(n3860), .Y(n2747) );
  OAI222XL U3622 ( .A0(n1384), .A1(n4009), .B0(n4047), .B1(n4006), .C0(n4301), 
        .C1(n3860), .Y(n2746) );
  OAI222XL U3623 ( .A0(n1385), .A1(n4009), .B0(n4049), .B1(n4006), .C0(n4300), 
        .C1(n3861), .Y(n2745) );
  OAI222XL U3624 ( .A0(n1386), .A1(n4009), .B0(n4051), .B1(n4006), .C0(n4299), 
        .C1(n3861), .Y(n2744) );
  OAI222XL U3625 ( .A0(n1387), .A1(n4009), .B0(n4053), .B1(n4006), .C0(n4298), 
        .C1(n3860), .Y(n2743) );
  OAI222XL U3626 ( .A0(n1388), .A1(n4009), .B0(n4055), .B1(n4006), .C0(n4297), 
        .C1(n3860), .Y(n2742) );
  OAI222XL U3627 ( .A0(n1389), .A1(n4009), .B0(n4057), .B1(n4006), .C0(n4296), 
        .C1(n3861), .Y(n2741) );
  OAI222XL U3628 ( .A0(n1390), .A1(n4009), .B0(n4059), .B1(n4006), .C0(n4295), 
        .C1(n3861), .Y(n2740) );
  OAI222XL U3629 ( .A0(n1391), .A1(n4009), .B0(n4062), .B1(n4008), .C0(n4294), 
        .C1(n3861), .Y(n2739) );
  OAI222XL U3630 ( .A0(n1392), .A1(n4009), .B0(n4065), .B1(n4008), .C0(n4293), 
        .C1(n3861), .Y(n2738) );
  OAI222XL U3631 ( .A0(n1393), .A1(n4009), .B0(n4068), .B1(n4008), .C0(n4292), 
        .C1(n3861), .Y(n2737) );
  OAI222XL U3632 ( .A0(n1394), .A1(n4009), .B0(n4071), .B1(n4008), .C0(n4291), 
        .C1(n3861), .Y(n2736) );
  OAI222XL U3633 ( .A0(n1395), .A1(n4009), .B0(n4074), .B1(n4008), .C0(n4290), 
        .C1(n3861), .Y(n2735) );
  OAI222XL U3634 ( .A0(n1396), .A1(n4009), .B0(n4077), .B1(n4008), .C0(n4289), 
        .C1(n3861), .Y(n2734) );
  OAI222XL U3635 ( .A0(n1397), .A1(n4010), .B0(n4080), .B1(n4008), .C0(n4288), 
        .C1(n3861), .Y(n2733) );
  OAI222XL U3636 ( .A0(n1398), .A1(n4010), .B0(n4083), .B1(n4008), .C0(n4287), 
        .C1(n3861), .Y(n2732) );
  OAI222XL U3637 ( .A0(n1399), .A1(n4010), .B0(n4086), .B1(n4008), .C0(n4286), 
        .C1(n3861), .Y(n2731) );
  OAI222XL U3638 ( .A0(n1400), .A1(n4010), .B0(n4089), .B1(n4008), .C0(n4285), 
        .C1(n3861), .Y(n2730) );
  OAI222XL U3639 ( .A0(n1401), .A1(n4010), .B0(n4092), .B1(n4008), .C0(n4284), 
        .C1(n3864), .Y(n2729) );
  OAI222XL U3640 ( .A0(n1402), .A1(n4010), .B0(n4095), .B1(n4008), .C0(n4283), 
        .C1(n3861), .Y(n2728) );
  OAI222XL U3641 ( .A0(n1403), .A1(n4010), .B0(n4098), .B1(n4007), .C0(n4282), 
        .C1(n3861), .Y(n2727) );
  OAI222XL U3642 ( .A0(n1404), .A1(n4010), .B0(n4101), .B1(n4007), .C0(n4281), 
        .C1(n3858), .Y(n2726) );
  OAI222XL U3643 ( .A0(n1405), .A1(n4010), .B0(n4104), .B1(n4007), .C0(n4280), 
        .C1(n3862), .Y(n2725) );
  OAI222XL U3644 ( .A0(n1406), .A1(n4010), .B0(n4107), .B1(n4007), .C0(n4279), 
        .C1(n3865), .Y(n2724) );
  OAI222XL U3645 ( .A0(n1407), .A1(n4010), .B0(n4110), .B1(n4007), .C0(n4278), 
        .C1(n3863), .Y(n2723) );
  OAI222XL U3646 ( .A0(n1408), .A1(n4010), .B0(n4029), .B1(n4007), .C0(n4277), 
        .C1(n3861), .Y(n2722) );
  OAI222XL U3647 ( .A0(n1409), .A1(n4010), .B0(n4031), .B1(n4007), .C0(n4276), 
        .C1(n3858), .Y(n2721) );
  OAI222XL U3648 ( .A0(n1410), .A1(n4010), .B0(n4033), .B1(n4007), .C0(n4275), 
        .C1(n3865), .Y(n2720) );
  OAI222XL U3649 ( .A0(n1411), .A1(n4010), .B0(n4035), .B1(n4007), .C0(n4274), 
        .C1(n3859), .Y(n2719) );
  OAI222XL U3650 ( .A0(n1412), .A1(n4010), .B0(n4037), .B1(n4007), .C0(n4273), 
        .C1(n3863), .Y(n2718) );
  OAI222XL U3651 ( .A0(n1413), .A1(n4009), .B0(n4039), .B1(n4007), .C0(n4272), 
        .C1(n3859), .Y(n2717) );
  OAI222XL U3652 ( .A0(n1414), .A1(n195), .B0(n4041), .B1(n4007), .C0(n4271), 
        .C1(n3864), .Y(n2716) );
  OAI222XL U3653 ( .A0(n1511), .A1(n4020), .B0(n4044), .B1(n4017), .C0(n4302), 
        .C1(n3872), .Y(n2619) );
  OAI222XL U3654 ( .A0(n1512), .A1(n4020), .B0(n4047), .B1(n4017), .C0(n4301), 
        .C1(n3873), .Y(n2618) );
  OAI222XL U3655 ( .A0(n1513), .A1(n4020), .B0(n4049), .B1(n4017), .C0(n4300), 
        .C1(n3872), .Y(n2617) );
  OAI222XL U3656 ( .A0(n1514), .A1(n4020), .B0(n4051), .B1(n4017), .C0(n4299), 
        .C1(n3872), .Y(n2616) );
  OAI222XL U3657 ( .A0(n1515), .A1(n4020), .B0(n4053), .B1(n4017), .C0(n4298), 
        .C1(n3873), .Y(n2615) );
  OAI222XL U3658 ( .A0(n1516), .A1(n4020), .B0(n4055), .B1(n4017), .C0(n4297), 
        .C1(n3873), .Y(n2614) );
  OAI222XL U3659 ( .A0(n1517), .A1(n4020), .B0(n4057), .B1(n4017), .C0(n4296), 
        .C1(n3872), .Y(n2613) );
  OAI222XL U3660 ( .A0(n1518), .A1(n4020), .B0(n4059), .B1(n4017), .C0(n4295), 
        .C1(n3873), .Y(n2612) );
  OAI222XL U3661 ( .A0(n1519), .A1(n4020), .B0(n4062), .B1(n4019), .C0(n4294), 
        .C1(n3873), .Y(n2611) );
  OAI222XL U3662 ( .A0(n1520), .A1(n4020), .B0(n4065), .B1(n4019), .C0(n4293), 
        .C1(n3873), .Y(n2610) );
  OAI222XL U3663 ( .A0(n1521), .A1(n4020), .B0(n4068), .B1(n4019), .C0(n4292), 
        .C1(n3873), .Y(n2609) );
  OAI222XL U3664 ( .A0(n1522), .A1(n4020), .B0(n4071), .B1(n4019), .C0(n4291), 
        .C1(n3873), .Y(n2608) );
  OAI222XL U3665 ( .A0(n1523), .A1(n4020), .B0(n4074), .B1(n4019), .C0(n4290), 
        .C1(n3873), .Y(n2607) );
  OAI222XL U3666 ( .A0(n1524), .A1(n4020), .B0(n4077), .B1(n4019), .C0(n4289), 
        .C1(n3873), .Y(n2606) );
  OAI222XL U3667 ( .A0(n1525), .A1(n4021), .B0(n4080), .B1(n4019), .C0(n4288), 
        .C1(n3873), .Y(n2605) );
  OAI222XL U3668 ( .A0(n1526), .A1(n4021), .B0(n4083), .B1(n4019), .C0(n4287), 
        .C1(n3873), .Y(n2604) );
  OAI222XL U3669 ( .A0(n1527), .A1(n4021), .B0(n4086), .B1(n4019), .C0(n4286), 
        .C1(n3873), .Y(n2603) );
  OAI222XL U3670 ( .A0(n1528), .A1(n4021), .B0(n4089), .B1(n4019), .C0(n4285), 
        .C1(n3873), .Y(n2602) );
  OAI222XL U3671 ( .A0(n1529), .A1(n4021), .B0(n4092), .B1(n4019), .C0(n4284), 
        .C1(n3874), .Y(n2601) );
  OAI222XL U3672 ( .A0(n1530), .A1(n4021), .B0(n4095), .B1(n4019), .C0(n4283), 
        .C1(n3873), .Y(n2600) );
  OAI222XL U3673 ( .A0(n1531), .A1(n4021), .B0(n4098), .B1(n4018), .C0(n4282), 
        .C1(n3874), .Y(n2599) );
  OAI222XL U3674 ( .A0(n1532), .A1(n4021), .B0(n4101), .B1(n4018), .C0(n4281), 
        .C1(n3874), .Y(n2598) );
  OAI222XL U3675 ( .A0(n1533), .A1(n4021), .B0(n4104), .B1(n4018), .C0(n4280), 
        .C1(n3873), .Y(n2597) );
  OAI222XL U3676 ( .A0(n1534), .A1(n4021), .B0(n4107), .B1(n4018), .C0(n4279), 
        .C1(n3874), .Y(n2596) );
  OAI222XL U3677 ( .A0(n1535), .A1(n4021), .B0(n4110), .B1(n4018), .C0(n4278), 
        .C1(n3874), .Y(n2595) );
  OAI222XL U3678 ( .A0(n1536), .A1(n4021), .B0(n3214), .B1(n4018), .C0(n4277), 
        .C1(n3874), .Y(n2594) );
  OAI222XL U3679 ( .A0(n1537), .A1(n4021), .B0(n3215), .B1(n4018), .C0(n4276), 
        .C1(n3874), .Y(n2593) );
  OAI222XL U3680 ( .A0(n1538), .A1(n4021), .B0(n3216), .B1(n4018), .C0(n4275), 
        .C1(n3874), .Y(n2592) );
  OAI222XL U3681 ( .A0(n1539), .A1(n4021), .B0(n3205), .B1(n4018), .C0(n4274), 
        .C1(n3874), .Y(n2591) );
  OAI222XL U3682 ( .A0(n1540), .A1(n4021), .B0(n3206), .B1(n4018), .C0(n4273), 
        .C1(n3874), .Y(n2590) );
  OAI222XL U3683 ( .A0(n1541), .A1(n4021), .B0(n3207), .B1(n4018), .C0(n4272), 
        .C1(n3874), .Y(n2589) );
  OAI222XL U3684 ( .A0(n1542), .A1(n4021), .B0(n3208), .B1(n4018), .C0(n4271), 
        .C1(n3874), .Y(n2588) );
  OAI222XL U3685 ( .A0(n1639), .A1(n4042), .B0(n4044), .B1(n3173), .C0(n3888), 
        .C1(n4302), .Y(n2491) );
  OAI222XL U3686 ( .A0(n1640), .A1(n4042), .B0(n4047), .B1(n3173), .C0(n3888), 
        .C1(n4301), .Y(n2490) );
  OAI222XL U3687 ( .A0(n1641), .A1(n4042), .B0(n4049), .B1(n3173), .C0(n3888), 
        .C1(n4300), .Y(n2489) );
  OAI222XL U3688 ( .A0(n1642), .A1(n4042), .B0(n4051), .B1(n3173), .C0(n3888), 
        .C1(n4299), .Y(n2488) );
  OAI222XL U3689 ( .A0(n1643), .A1(n4042), .B0(n4053), .B1(n3173), .C0(n3888), 
        .C1(n4298), .Y(n2487) );
  OAI222XL U3690 ( .A0(n1644), .A1(n4042), .B0(n4055), .B1(n3173), .C0(n3888), 
        .C1(n4297), .Y(n2486) );
  OAI222XL U3691 ( .A0(n1645), .A1(n4042), .B0(n4057), .B1(n3173), .C0(n3888), 
        .C1(n4296), .Y(n2485) );
  OAI222XL U3692 ( .A0(n1646), .A1(n4042), .B0(n4059), .B1(n3173), .C0(n3888), 
        .C1(n4295), .Y(n2484) );
  OAI222XL U3693 ( .A0(n1647), .A1(n4042), .B0(n4062), .B1(n3173), .C0(n3888), 
        .C1(n4294), .Y(n2483) );
  OAI222XL U3694 ( .A0(n1648), .A1(n4042), .B0(n4065), .B1(n3173), .C0(n3888), 
        .C1(n4293), .Y(n2482) );
  OAI222XL U3695 ( .A0(n1649), .A1(n4042), .B0(n4068), .B1(n3173), .C0(n3888), 
        .C1(n4292), .Y(n2481) );
  OAI222XL U3696 ( .A0(n1650), .A1(n4042), .B0(n4071), .B1(n3173), .C0(n3888), 
        .C1(n4291), .Y(n2480) );
  OAI222XL U3697 ( .A0(n1651), .A1(n4042), .B0(n4074), .B1(n3173), .C0(n3889), 
        .C1(n4290), .Y(n2479) );
  OAI222XL U3698 ( .A0(n1652), .A1(n4042), .B0(n4077), .B1(n3173), .C0(n3889), 
        .C1(n4289), .Y(n2478) );
  OAI222XL U3699 ( .A0(n1653), .A1(n4042), .B0(n4080), .B1(n3173), .C0(n3889), 
        .C1(n4288), .Y(n2477) );
  OAI222XL U3700 ( .A0(n1654), .A1(n4042), .B0(n4083), .B1(n3173), .C0(n3889), 
        .C1(n4287), .Y(n2476) );
  OAI222XL U3701 ( .A0(n1655), .A1(n4042), .B0(n4086), .B1(n3173), .C0(n3889), 
        .C1(n4286), .Y(n2475) );
  OAI222XL U3702 ( .A0(n1656), .A1(n4042), .B0(n4089), .B1(n3173), .C0(n3889), 
        .C1(n4285), .Y(n2474) );
  OAI222XL U3703 ( .A0(n1657), .A1(n4042), .B0(n4092), .B1(n3173), .C0(n3889), 
        .C1(n4284), .Y(n2473) );
  OAI222XL U3704 ( .A0(n1658), .A1(n4042), .B0(n4095), .B1(n3173), .C0(n3889), 
        .C1(n4283), .Y(n2472) );
  OAI222XL U3705 ( .A0(n1659), .A1(n4042), .B0(n4098), .B1(n3173), .C0(n3889), 
        .C1(n4282), .Y(n2471) );
  OAI222XL U3706 ( .A0(n1660), .A1(n4042), .B0(n4101), .B1(n3173), .C0(n3889), 
        .C1(n4281), .Y(n2470) );
  OAI222XL U3707 ( .A0(n1661), .A1(n4042), .B0(n4104), .B1(n3173), .C0(n3889), 
        .C1(n4280), .Y(n2469) );
  OAI222XL U3708 ( .A0(n1662), .A1(n4042), .B0(n4107), .B1(n3173), .C0(n3889), 
        .C1(n4279), .Y(n2468) );
  OAI222XL U3709 ( .A0(n1663), .A1(n4042), .B0(n4110), .B1(n3173), .C0(n3889), 
        .C1(n4278), .Y(n2467) );
  OAI222XL U3710 ( .A0(n1664), .A1(n4042), .B0(n3173), .B1(n4028), .C0(n3889), 
        .C1(n4277), .Y(n2466) );
  OAI222XL U3711 ( .A0(n1665), .A1(n4042), .B0(n3173), .B1(n4030), .C0(n3889), 
        .C1(n4276), .Y(n2465) );
  OAI222XL U3712 ( .A0(n1666), .A1(n4042), .B0(n3173), .B1(n4032), .C0(n3889), 
        .C1(n4275), .Y(n2464) );
  OAI222XL U3713 ( .A0(n1667), .A1(n4042), .B0(n3173), .B1(n4034), .C0(n3890), 
        .C1(n4274), .Y(n2463) );
  OAI222XL U3714 ( .A0(n1668), .A1(n4042), .B0(n3173), .B1(n4036), .C0(n3890), 
        .C1(n4273), .Y(n2462) );
  OAI222XL U3715 ( .A0(n1669), .A1(n4042), .B0(n3173), .B1(n4038), .C0(n3890), 
        .C1(n4272), .Y(n2461) );
  OAI222XL U3716 ( .A0(n1670), .A1(n4042), .B0(n3173), .B1(n4040), .C0(n3890), 
        .C1(n4271), .Y(n2460) );
  MXI2X1 U3717 ( .A(n3324), .B(n3325), .S0(n3658), .Y(N224) );
  MXI2X1 U3718 ( .A(n3306), .B(n3307), .S0(n3657), .Y(N215) );
  MXI4X1 U3719 ( .A(\tag[0][16] ), .B(\tag[1][16] ), .C(\tag[2][16] ), .D(
        \tag[3][16] ), .S0(n3275), .S1(n3631), .Y(n3306) );
  MXI4X1 U3720 ( .A(\tag[4][16] ), .B(\tag[5][16] ), .C(\tag[6][16] ), .D(
        \tag[7][16] ), .S0(n3275), .S1(n3631), .Y(n3307) );
  MXI2X1 U3721 ( .A(n3298), .B(n3299), .S0(n3657), .Y(N210) );
  MXI4X1 U3722 ( .A(\tag[4][21] ), .B(\tag[5][21] ), .C(\tag[6][21] ), .D(
        \tag[7][21] ), .S0(n3602), .S1(n3631), .Y(n3299) );
  MXI4X1 U3723 ( .A(\tag[0][21] ), .B(\tag[1][21] ), .C(\tag[2][21] ), .D(
        \tag[3][21] ), .S0(n3275), .S1(n3631), .Y(n3298) );
  MXI2X1 U3724 ( .A(n3296), .B(n3297), .S0(n3657), .Y(N209) );
  MXI4X1 U3725 ( .A(\tag[0][22] ), .B(\tag[1][22] ), .C(\tag[2][22] ), .D(
        \tag[3][22] ), .S0(n3602), .S1(n3630), .Y(n3296) );
  MXI4X1 U3726 ( .A(\tag[4][22] ), .B(\tag[5][22] ), .C(\tag[6][22] ), .D(
        \tag[7][22] ), .S0(n3602), .S1(n3630), .Y(n3297) );
  MXI2X1 U3727 ( .A(n3294), .B(n3295), .S0(n3657), .Y(N208) );
  MXI4X1 U3728 ( .A(\tag[0][23] ), .B(\tag[1][23] ), .C(\tag[2][23] ), .D(
        \tag[3][23] ), .S0(n3602), .S1(n3630), .Y(n3294) );
  MXI4X1 U3729 ( .A(\tag[4][23] ), .B(\tag[5][23] ), .C(\tag[6][23] ), .D(
        \tag[7][23] ), .S0(n3602), .S1(n3630), .Y(n3295) );
  MXI2X1 U3730 ( .A(n3328), .B(n3329), .S0(n3658), .Y(N226) );
  MXI4X1 U3731 ( .A(\tag[0][24] ), .B(\tag[1][24] ), .C(\tag[2][24] ), .D(
        \tag[3][24] ), .S0(n3602), .S1(n3630), .Y(n3292) );
  MXI4X1 U3732 ( .A(\tag[4][24] ), .B(\tag[5][24] ), .C(\tag[6][24] ), .D(
        \tag[7][24] ), .S0(n3602), .S1(n3630), .Y(n3293) );
  MXI2X1 U3733 ( .A(n3302), .B(n3303), .S0(n3657), .Y(N213) );
  MXI4X1 U3734 ( .A(\tag[0][18] ), .B(\tag[1][18] ), .C(\tag[2][18] ), .D(
        \tag[3][18] ), .S0(n3275), .S1(n3631), .Y(n3302) );
  MXI4X1 U3735 ( .A(\tag[4][18] ), .B(\tag[5][18] ), .C(\tag[6][18] ), .D(
        \tag[7][18] ), .S0(n3275), .S1(n3631), .Y(n3303) );
  MXI2X1 U3736 ( .A(n3326), .B(n3327), .S0(n3658), .Y(N225) );
  MXI2X1 U3737 ( .A(n3334), .B(n3335), .S0(n3659), .Y(N229) );
  MXI2X1 U3738 ( .A(n3330), .B(n3331), .S0(n3658), .Y(N227) );
  MXI2X1 U3739 ( .A(n3322), .B(n3323), .S0(n3658), .Y(N223) );
  MXI4X1 U3740 ( .A(\tag[0][8] ), .B(\tag[1][8] ), .C(\tag[2][8] ), .D(
        \tag[3][8] ), .S0(n3605), .S1(n3633), .Y(n3322) );
  MXI4X1 U3741 ( .A(\tag[4][8] ), .B(\tag[5][8] ), .C(\tag[6][8] ), .D(
        \tag[7][8] ), .S0(n3605), .S1(n3633), .Y(n3323) );
  MXI2X1 U3742 ( .A(n3314), .B(n3315), .S0(n3658), .Y(N219) );
  MXI4X1 U3743 ( .A(\tag[0][12] ), .B(\tag[1][12] ), .C(\tag[2][12] ), .D(
        \tag[3][12] ), .S0(n3605), .S1(n3632), .Y(n3314) );
  MXI4X1 U3744 ( .A(\tag[4][12] ), .B(\tag[5][12] ), .C(\tag[6][12] ), .D(
        \tag[7][12] ), .S0(n3605), .S1(n3632), .Y(n3315) );
  MXI2X1 U3745 ( .A(n3332), .B(n3333), .S0(n3659), .Y(N228) );
  MXI4X1 U3746 ( .A(\tag[0][3] ), .B(\tag[1][3] ), .C(\tag[2][3] ), .D(
        \tag[3][3] ), .S0(n3605), .S1(n3634), .Y(n3332) );
  MXI4X1 U3747 ( .A(\tag[4][3] ), .B(\tag[5][3] ), .C(\tag[6][3] ), .D(
        \tag[7][3] ), .S0(n3605), .S1(n3634), .Y(n3333) );
  MXI2X1 U3748 ( .A(n3300), .B(n3301), .S0(n3657), .Y(N212) );
  MXI2X1 U3749 ( .A(n3320), .B(n3321), .S0(n3658), .Y(N222) );
  MXI4X1 U3750 ( .A(\tag[0][9] ), .B(\tag[1][9] ), .C(\tag[2][9] ), .D(
        \tag[3][9] ), .S0(n3605), .S1(n3633), .Y(n3320) );
  MXI4X1 U3751 ( .A(\tag[4][9] ), .B(\tag[5][9] ), .C(\tag[6][9] ), .D(
        \tag[7][9] ), .S0(n3605), .S1(n3633), .Y(n3321) );
  MXI4X1 U3752 ( .A(\tag[4][15] ), .B(\tag[5][15] ), .C(\tag[6][15] ), .D(
        \tag[7][15] ), .S0(n3603), .S1(n3632), .Y(n3309) );
  MXI2X1 U3753 ( .A(n3310), .B(n3311), .S0(n3658), .Y(N217) );
  MXI4X1 U3754 ( .A(\tag[0][14] ), .B(\tag[1][14] ), .C(\tag[2][14] ), .D(
        \tag[3][14] ), .S0(n3604), .S1(n3632), .Y(n3310) );
  MXI4X1 U3755 ( .A(\tag[4][14] ), .B(\tag[5][14] ), .C(\tag[6][14] ), .D(
        \tag[7][14] ), .S0(n3604), .S1(n3632), .Y(n3311) );
  MXI2X1 U3756 ( .A(n3312), .B(n3313), .S0(n3658), .Y(N218) );
  MXI4X1 U3757 ( .A(\tag[0][13] ), .B(\tag[1][13] ), .C(\tag[2][13] ), .D(
        \tag[3][13] ), .S0(n3604), .S1(n3632), .Y(n3312) );
  MXI4X1 U3758 ( .A(\tag[4][13] ), .B(\tag[5][13] ), .C(\tag[6][13] ), .D(
        \tag[7][13] ), .S0(n3604), .S1(n3632), .Y(n3313) );
  MXI2X1 U3759 ( .A(n3318), .B(n3319), .S0(n3658), .Y(N221) );
  MXI4X1 U3760 ( .A(\tag[0][10] ), .B(\tag[1][10] ), .C(\tag[2][10] ), .D(
        \tag[3][10] ), .S0(n3604), .S1(n3632), .Y(n3318) );
  MXI4X1 U3761 ( .A(\tag[4][10] ), .B(\tag[5][10] ), .C(\tag[6][10] ), .D(
        \tag[7][10] ), .S0(n3604), .S1(n3632), .Y(n3319) );
  MXI2X1 U3762 ( .A(n3316), .B(n3317), .S0(n3658), .Y(N220) );
  MXI4X1 U3763 ( .A(\tag[0][11] ), .B(\tag[1][11] ), .C(\tag[2][11] ), .D(
        \tag[3][11] ), .S0(n3604), .S1(n3632), .Y(n3316) );
  MXI4X1 U3764 ( .A(\tag[4][11] ), .B(\tag[5][11] ), .C(\tag[6][11] ), .D(
        \tag[7][11] ), .S0(n3604), .S1(n3632), .Y(n3317) );
  MXI2X1 U3765 ( .A(n3338), .B(n3339), .S0(n3659), .Y(N231) );
  MXI4X1 U3766 ( .A(\tag[0][0] ), .B(\tag[1][0] ), .C(\tag[2][0] ), .D(
        \tag[3][0] ), .S0(n3606), .S1(n3634), .Y(n3338) );
  MXI4X1 U3767 ( .A(\tag[4][0] ), .B(\tag[5][0] ), .C(\tag[6][0] ), .D(
        \tag[7][0] ), .S0(n3606), .S1(n3634), .Y(n3339) );
  XNOR2X1 U3768 ( .A(N223), .B(proc_addr[13]), .Y(n385) );
  XNOR2X1 U3769 ( .A(N211), .B(proc_addr[25]), .Y(n384) );
  XNOR2X1 U3770 ( .A(N219), .B(proc_addr[17]), .Y(n383) );
  XNOR2X1 U3771 ( .A(N231), .B(proc_addr[5]), .Y(n378) );
  NAND4X1 U3772 ( .A(n376), .B(n377), .C(n378), .D(N232), .Y(n372) );
  MXI2X1 U3773 ( .A(n3290), .B(n3291), .S0(n3657), .Y(N232) );
  XNOR2X1 U3774 ( .A(N228), .B(proc_addr[8]), .Y(n376) );
  OAI222XL U3775 ( .A0(n3999), .A1(n4148), .B0(n4149), .B1(n3998), .C0(n1326), 
        .C1(n3805), .Y(n2837) );
  OAI222XL U3776 ( .A0(n3999), .A1(n4147), .B0(n3251), .B1(n3998), .C0(n1327), 
        .C1(n3805), .Y(n2836) );
  OAI222XL U3777 ( .A0(n3999), .A1(n4146), .B0(n4150), .B1(n3998), .C0(n1328), 
        .C1(n3805), .Y(n2835) );
  OAI222XL U3778 ( .A0(n3999), .A1(n4145), .B0(n4151), .B1(n3998), .C0(n1329), 
        .C1(n3805), .Y(n2834) );
  OAI222XL U3779 ( .A0(n3999), .A1(n4144), .B0(n4152), .B1(n208), .C0(n1330), 
        .C1(n3805), .Y(n2833) );
  OAI222XL U3780 ( .A0(n205), .A1(n4143), .B0(n4153), .B1(n208), .C0(n1331), 
        .C1(n3805), .Y(n2832) );
  OAI222XL U3781 ( .A0(n205), .A1(n4142), .B0(n4154), .B1(n208), .C0(n1332), 
        .C1(n3805), .Y(n2831) );
  OAI222XL U3782 ( .A0(n205), .A1(n4141), .B0(n4155), .B1(n208), .C0(n1333), 
        .C1(n3805), .Y(n2830) );
  OAI222XL U3783 ( .A0(n205), .A1(n4140), .B0(n4156), .B1(n208), .C0(n1334), 
        .C1(n3805), .Y(n2829) );
  OAI222XL U3784 ( .A0(n205), .A1(n4139), .B0(n4157), .B1(n208), .C0(n1335), 
        .C1(n3805), .Y(n2828) );
  OAI222XL U3785 ( .A0(n3999), .A1(n4138), .B0(n4158), .B1(n3998), .C0(n1336), 
        .C1(n3805), .Y(n2827) );
  OAI222XL U3786 ( .A0(n3999), .A1(n4137), .B0(n4159), .B1(n3998), .C0(n1337), 
        .C1(n3805), .Y(n2826) );
  OAI222XL U3787 ( .A0(n3999), .A1(n4136), .B0(n4160), .B1(n3998), .C0(n1338), 
        .C1(n3806), .Y(n2825) );
  OAI222XL U3788 ( .A0(n3999), .A1(n4135), .B0(n4161), .B1(n3998), .C0(n1339), 
        .C1(n3806), .Y(n2824) );
  OAI222XL U3789 ( .A0(n3999), .A1(n4134), .B0(n4162), .B1(n3998), .C0(n1340), 
        .C1(n3806), .Y(n2823) );
  OAI222XL U3790 ( .A0(n3999), .A1(n4133), .B0(n3248), .B1(n3998), .C0(n1341), 
        .C1(n3806), .Y(n2822) );
  OAI222XL U3791 ( .A0(n3999), .A1(n4132), .B0(n4163), .B1(n3998), .C0(n1342), 
        .C1(n3806), .Y(n2821) );
  OAI222XL U3792 ( .A0(n3999), .A1(n4131), .B0(n4164), .B1(n3998), .C0(n1343), 
        .C1(n3806), .Y(n2820) );
  OAI222XL U3793 ( .A0(n3999), .A1(n4130), .B0(n4165), .B1(n3998), .C0(n1344), 
        .C1(n3806), .Y(n2819) );
  OAI222XL U3794 ( .A0(n3999), .A1(n4129), .B0(n4166), .B1(n3998), .C0(n1345), 
        .C1(n3806), .Y(n2818) );
  OAI222XL U3795 ( .A0(n3999), .A1(n4128), .B0(n4167), .B1(n3998), .C0(n1346), 
        .C1(n3806), .Y(n2817) );
  OAI222XL U3796 ( .A0(n3999), .A1(n4127), .B0(n4168), .B1(n3998), .C0(n1347), 
        .C1(n3806), .Y(n2816) );
  OAI222XL U3797 ( .A0(n3999), .A1(n4126), .B0(n4169), .B1(n3998), .C0(n1348), 
        .C1(n3806), .Y(n2815) );
  OAI222XL U3798 ( .A0(n3999), .A1(n4125), .B0(n4170), .B1(n3998), .C0(n1349), 
        .C1(n3806), .Y(n2814) );
  OAI222XL U3799 ( .A0(n3999), .A1(n4124), .B0(n4171), .B1(n3998), .C0(n1350), 
        .C1(n3806), .Y(n2813) );
  OAI32X1 U3800 ( .A0(n268), .A1(n4172), .A2(n269), .B0(n1322), .B1(n270), .Y(
        n2969) );
  NAND3X1 U3801 ( .A(n4303), .B(n3667), .C(n270), .Y(n268) );
  NOR2X1 U3802 ( .A(n4306), .B(state[0]), .Y(n288) );
  NOR2X1 U3803 ( .A(state[1]), .B(state[0]), .Y(n303) );
  AOI211X1 U3804 ( .A0(n286), .A1(n287), .B0(n288), .C0(n289), .Y(n3170) );
  OR2X1 U3805 ( .A(n290), .B(mem_ready), .Y(n286) );
  OAI21XL U3806 ( .A0(N233), .A1(n269), .B0(n290), .Y(n287) );
  OAI22XL U3807 ( .A0(n1323), .A1(n3805), .B0(n261), .B1(n4119), .Y(n2840) );
  OAI22XL U3808 ( .A0(n1324), .A1(n3805), .B0(n261), .B1(n4117), .Y(n2839) );
  OAI22XL U3809 ( .A0(n1325), .A1(n3805), .B0(n261), .B1(n4115), .Y(n2838) );
  OAI2BB2XL U3810 ( .B0(n301), .B1(n1120), .A0N(n3280), .A1N(n301), .Y(n1715)
         );
  NAND4X1 U3811 ( .A(n269), .B(n3667), .C(n4303), .D(n302), .Y(n3280) );
  NAND2X1 U3812 ( .A(n4121), .B(n302), .Y(n301) );
  OAI22XL U3813 ( .A0(n190), .A1(n306), .B0(n1112), .B1(n319), .Y(n1723) );
  NOR2X1 U3814 ( .A(n3668), .B(n190), .Y(n319) );
  OAI22XL U3815 ( .A0(n139), .A1(n306), .B0(n1113), .B1(n318), .Y(n1722) );
  NOR2X1 U3816 ( .A(n3668), .B(n139), .Y(n318) );
  OAI22XL U3817 ( .A0(n101), .A1(n306), .B0(n1114), .B1(n317), .Y(n1721) );
  NOR2X1 U3818 ( .A(n3668), .B(n101), .Y(n317) );
  OAI22XL U3819 ( .A0(n315), .A1(n306), .B0(n1115), .B1(n316), .Y(n1720) );
  NOR2X1 U3820 ( .A(n3668), .B(n315), .Y(n316) );
  OAI22XL U3821 ( .A0(n313), .A1(n306), .B0(n1116), .B1(n314), .Y(n1719) );
  NOR2X1 U3822 ( .A(n3668), .B(n313), .Y(n314) );
  OAI22XL U3823 ( .A0(n311), .A1(n306), .B0(n1117), .B1(n312), .Y(n1718) );
  NOR2X1 U3824 ( .A(n3668), .B(n311), .Y(n312) );
  OAI22XL U3825 ( .A0(n309), .A1(n306), .B0(n1118), .B1(n310), .Y(n1717) );
  NOR2X1 U3826 ( .A(n3668), .B(n309), .Y(n310) );
  OAI22XL U3827 ( .A0(n305), .A1(n306), .B0(n1119), .B1(n307), .Y(n1716) );
  NOR2X1 U3828 ( .A(n3668), .B(n305), .Y(n307) );
  OAI2BB2XL U3829 ( .B0(n4307), .B1(n202), .A0N(n202), .A1N(proc_write), .Y(
        n2780) );
  OAI2BB2XL U3830 ( .B0(n4004), .B1(n1374), .A0N(N183), .A1N(n4004), .Y(n2756)
         );
  MX4X1 U3831 ( .A(N151), .B(N119), .C(N87), .D(N55), .S0(n3286), .S1(n3288), 
        .Y(N183) );
  OAI2BB2XL U3832 ( .B0(n4004), .B1(n1376), .A0N(N181), .A1N(n4005), .Y(n2754)
         );
  MX4X1 U3833 ( .A(N149), .B(N117), .C(N85), .D(N53), .S0(n3287), .S1(n3289), 
        .Y(N181) );
  OAI2BB2XL U3834 ( .B0(n4004), .B1(n1377), .A0N(N180), .A1N(n4005), .Y(n2753)
         );
  MX4X1 U3835 ( .A(N148), .B(N116), .C(N84), .D(N52), .S0(n3286), .S1(n3288), 
        .Y(N180) );
  OAI2BB2XL U3836 ( .B0(n4004), .B1(n1378), .A0N(N179), .A1N(n4005), .Y(n2752)
         );
  MX4X1 U3837 ( .A(N147), .B(N115), .C(N83), .D(N51), .S0(n3285), .S1(n3289), 
        .Y(N179) );
  OAI2BB2XL U3838 ( .B0(n4004), .B1(n1379), .A0N(N178), .A1N(n4005), .Y(n2751)
         );
  MX4X1 U3839 ( .A(N146), .B(N114), .C(N82), .D(N50), .S0(n3285), .S1(n3288), 
        .Y(N178) );
  OAI2BB2XL U3840 ( .B0(n4004), .B1(n1380), .A0N(N177), .A1N(n4005), .Y(n2750)
         );
  MX4X1 U3841 ( .A(N145), .B(N113), .C(N81), .D(N49), .S0(n3285), .S1(n3289), 
        .Y(N177) );
  OAI2BB2XL U3842 ( .B0(n4004), .B1(n1381), .A0N(N176), .A1N(n4003), .Y(n2749)
         );
  MX4X1 U3843 ( .A(N144), .B(N112), .C(N80), .D(N48), .S0(N45), .S1(n3288), 
        .Y(N176) );
  OAI2BB2XL U3844 ( .B0(n4004), .B1(n1382), .A0N(N175), .A1N(n4005), .Y(n2748)
         );
  MX4X1 U3845 ( .A(N143), .B(N111), .C(N79), .D(N47), .S0(N45), .S1(n3289), 
        .Y(N175) );
  OAI2BB2XL U3846 ( .B0(n4004), .B1(n1351), .A0N(N206), .A1N(n4003), .Y(n2779)
         );
  MX4X1 U3847 ( .A(N174), .B(N142), .C(N110), .D(N78), .S0(n3287), .S1(n3289), 
        .Y(N206) );
  OAI2BB2XL U3848 ( .B0(n4003), .B1(n1352), .A0N(N205), .A1N(n4005), .Y(n2778)
         );
  MX4X1 U3849 ( .A(N173), .B(N141), .C(N109), .D(N77), .S0(n3287), .S1(n3289), 
        .Y(N205) );
  OAI2BB2XL U3850 ( .B0(n4003), .B1(n1353), .A0N(N204), .A1N(n4003), .Y(n2777)
         );
  MX4X1 U3851 ( .A(N172), .B(N140), .C(N108), .D(N76), .S0(n3287), .S1(n3289), 
        .Y(N204) );
  OAI2BB2XL U3852 ( .B0(n4003), .B1(n1354), .A0N(N203), .A1N(n4005), .Y(n2776)
         );
  MX4X1 U3853 ( .A(N171), .B(N139), .C(N107), .D(N75), .S0(n3287), .S1(n3289), 
        .Y(N203) );
  OAI2BB2XL U3854 ( .B0(n4003), .B1(n1355), .A0N(N202), .A1N(n4005), .Y(n2775)
         );
  MX4X1 U3855 ( .A(N170), .B(N138), .C(N106), .D(N74), .S0(n3287), .S1(n3289), 
        .Y(N202) );
  OAI2BB2XL U3856 ( .B0(n4003), .B1(n1356), .A0N(N201), .A1N(n4005), .Y(n2774)
         );
  MX4X1 U3857 ( .A(N169), .B(N137), .C(N105), .D(N73), .S0(n3287), .S1(n3289), 
        .Y(N201) );
  OAI2BB2XL U3858 ( .B0(n4003), .B1(n1357), .A0N(N200), .A1N(n4005), .Y(n2773)
         );
  MX4X1 U3859 ( .A(N168), .B(N136), .C(N104), .D(N72), .S0(n3287), .S1(n3289), 
        .Y(N200) );
  OAI2BB2XL U3860 ( .B0(n4003), .B1(n1358), .A0N(N199), .A1N(n4005), .Y(n2772)
         );
  MX4X1 U3861 ( .A(N167), .B(N135), .C(N103), .D(N71), .S0(n3287), .S1(n3289), 
        .Y(N199) );
  OAI2BB2XL U3862 ( .B0(n4003), .B1(n1359), .A0N(N198), .A1N(n4005), .Y(n2771)
         );
  MX4X1 U3863 ( .A(N166), .B(N134), .C(N102), .D(N70), .S0(n3287), .S1(n3289), 
        .Y(N198) );
  OAI2BB2XL U3864 ( .B0(n4003), .B1(n1360), .A0N(N197), .A1N(n4005), .Y(n2770)
         );
  MX4X1 U3865 ( .A(N165), .B(N133), .C(N101), .D(N69), .S0(n3287), .S1(n3289), 
        .Y(N197) );
  OAI2BB2XL U3866 ( .B0(n4003), .B1(n1361), .A0N(N196), .A1N(n4005), .Y(n2769)
         );
  MX4X1 U3867 ( .A(N164), .B(N132), .C(N100), .D(N68), .S0(n3287), .S1(n3289), 
        .Y(N196) );
  OAI2BB2XL U3868 ( .B0(n4003), .B1(n1362), .A0N(N195), .A1N(n4005), .Y(n2768)
         );
  MX4X1 U3869 ( .A(N163), .B(N131), .C(N99), .D(N67), .S0(n3287), .S1(n3289), 
        .Y(N195) );
  OAI2BB2XL U3870 ( .B0(n4003), .B1(n1363), .A0N(N194), .A1N(n4005), .Y(n2767)
         );
  MX4X1 U3871 ( .A(N162), .B(N130), .C(N98), .D(N66), .S0(n3286), .S1(n3288), 
        .Y(N194) );
  OAI2BB2XL U3872 ( .B0(n4003), .B1(n1364), .A0N(N193), .A1N(n4005), .Y(n2766)
         );
  MX4X1 U3873 ( .A(N161), .B(N129), .C(N97), .D(N65), .S0(n3286), .S1(n3288), 
        .Y(N193) );
  OAI2BB2XL U3874 ( .B0(n4004), .B1(n1365), .A0N(N192), .A1N(n4005), .Y(n2765)
         );
  MX4X1 U3875 ( .A(N160), .B(N128), .C(N96), .D(N64), .S0(n3286), .S1(n3288), 
        .Y(N192) );
  OAI2BB2XL U3876 ( .B0(n4003), .B1(n1366), .A0N(N191), .A1N(n4004), .Y(n2764)
         );
  MX4X1 U3877 ( .A(N159), .B(N127), .C(N95), .D(N63), .S0(n3286), .S1(n3288), 
        .Y(N191) );
  OAI2BB2XL U3878 ( .B0(n4004), .B1(n1367), .A0N(N190), .A1N(n4005), .Y(n2763)
         );
  MX4X1 U3879 ( .A(N158), .B(N126), .C(N94), .D(N62), .S0(n3286), .S1(n3288), 
        .Y(N190) );
  OAI2BB2XL U3880 ( .B0(n4003), .B1(n1368), .A0N(N189), .A1N(n4004), .Y(n2762)
         );
  MX4X1 U3881 ( .A(N157), .B(N125), .C(N93), .D(N61), .S0(n3286), .S1(n3288), 
        .Y(N189) );
  OAI2BB2XL U3882 ( .B0(n197), .B1(n1369), .A0N(N188), .A1N(n4004), .Y(n2761)
         );
  MX4X1 U3883 ( .A(N156), .B(N124), .C(N92), .D(N60), .S0(n3286), .S1(n3288), 
        .Y(N188) );
  OAI2BB2XL U3884 ( .B0(n197), .B1(n1370), .A0N(N187), .A1N(n4004), .Y(n2760)
         );
  MX4X1 U3885 ( .A(N155), .B(N123), .C(N91), .D(N59), .S0(n3286), .S1(n3288), 
        .Y(N187) );
  OAI2BB2XL U3886 ( .B0(n197), .B1(n1371), .A0N(N186), .A1N(n4004), .Y(n2759)
         );
  MX4X1 U3887 ( .A(N154), .B(N122), .C(N90), .D(N58), .S0(n3286), .S1(n3288), 
        .Y(N186) );
  OAI2BB2XL U3888 ( .B0(n197), .B1(n1372), .A0N(N185), .A1N(n4004), .Y(n2758)
         );
  MX4X1 U3889 ( .A(N153), .B(N121), .C(N89), .D(N57), .S0(n3286), .S1(n3288), 
        .Y(N185) );
  OAI2BB2XL U3890 ( .B0(n4004), .B1(n1373), .A0N(N184), .A1N(n4005), .Y(n2757)
         );
  MX4X1 U3891 ( .A(N152), .B(N120), .C(N88), .D(N56), .S0(n3286), .S1(n3288), 
        .Y(N184) );
  OAI2BB2XL U3892 ( .B0(n4003), .B1(n1375), .A0N(N182), .A1N(n4005), .Y(n2755)
         );
  MX4X1 U3893 ( .A(N150), .B(N118), .C(N86), .D(N54), .S0(N45), .S1(n3288), 
        .Y(N182) );
  NAND2X1 U3894 ( .A(mem_ready), .B(n288), .Y(n272) );
  OAI32X1 U3895 ( .A0(n297), .A1(n4304), .A2(n4121), .B0(n1121), .B1(n270), 
        .Y(n1714) );
  OA21XL U3896 ( .A0(N233), .A1(n269), .B0(n4303), .Y(n297) );
  AND3X2 U3897 ( .A(n3807), .B(n303), .C(proc_write), .Y(n3281) );
  INVX3 U3898 ( .A(proc_addr[7]), .Y(n4146) );
  INVX3 U3899 ( .A(proc_addr[9]), .Y(n4144) );
  INVX3 U3900 ( .A(proc_addr[10]), .Y(n4143) );
  INVX3 U3901 ( .A(proc_addr[11]), .Y(n4142) );
  INVX3 U3902 ( .A(proc_addr[12]), .Y(n4141) );
  INVX3 U3903 ( .A(proc_addr[21]), .Y(n4132) );
  INVX3 U3904 ( .A(proc_addr[22]), .Y(n4131) );
  INVX3 U3905 ( .A(proc_addr[23]), .Y(n4130) );
  INVX3 U3906 ( .A(proc_addr[26]), .Y(n4127) );
  INVX3 U3907 ( .A(proc_addr[27]), .Y(n4126) );
  INVX3 U3908 ( .A(proc_addr[28]), .Y(n4125) );
  INVX3 U3909 ( .A(proc_addr[29]), .Y(n4124) );
  AO22X1 U3910 ( .A0(N174), .A1(n3968), .B0(n3991), .B1(mem_wdata[0]), .Y(
        n2968) );
  AO22X1 U3911 ( .A0(N173), .A1(n3968), .B0(n3991), .B1(mem_wdata[1]), .Y(
        n2967) );
  AO22X1 U3912 ( .A0(N172), .A1(n3968), .B0(n3991), .B1(mem_wdata[2]), .Y(
        n2966) );
  AO22X1 U3913 ( .A0(N171), .A1(n3968), .B0(n3990), .B1(mem_wdata[3]), .Y(
        n2965) );
  AO22X1 U3914 ( .A0(N170), .A1(n3968), .B0(n3990), .B1(mem_wdata[4]), .Y(
        n2964) );
  AO22X1 U3915 ( .A0(N169), .A1(n3968), .B0(n3990), .B1(mem_wdata[5]), .Y(
        n2963) );
  AO22X1 U3916 ( .A0(N168), .A1(n3968), .B0(n3990), .B1(mem_wdata[6]), .Y(
        n2962) );
  AO22X1 U3917 ( .A0(N167), .A1(n3968), .B0(n3990), .B1(mem_wdata[7]), .Y(
        n2961) );
  AO22X1 U3918 ( .A0(N166), .A1(n3967), .B0(n3990), .B1(mem_wdata[8]), .Y(
        n2960) );
  AO22X1 U3919 ( .A0(N165), .A1(n3967), .B0(n3989), .B1(mem_wdata[9]), .Y(
        n2959) );
  AO22X1 U3920 ( .A0(N164), .A1(n3967), .B0(n3989), .B1(mem_wdata[10]), .Y(
        n2958) );
  AO22X1 U3921 ( .A0(N163), .A1(n3967), .B0(n3989), .B1(mem_wdata[11]), .Y(
        n2957) );
  AO22X1 U3922 ( .A0(N162), .A1(n3967), .B0(n3989), .B1(mem_wdata[12]), .Y(
        n2956) );
  AO22X1 U3923 ( .A0(N161), .A1(n3967), .B0(n3989), .B1(mem_wdata[13]), .Y(
        n2955) );
  AO22X1 U3924 ( .A0(N160), .A1(n3967), .B0(n3989), .B1(mem_wdata[14]), .Y(
        n2954) );
  AO22X1 U3925 ( .A0(N159), .A1(n3967), .B0(n3988), .B1(mem_wdata[15]), .Y(
        n2953) );
  AO22X1 U3926 ( .A0(N158), .A1(n3967), .B0(n3988), .B1(mem_wdata[16]), .Y(
        n2952) );
  AO22X1 U3927 ( .A0(N157), .A1(n3967), .B0(n3988), .B1(mem_wdata[17]), .Y(
        n2951) );
  AO22X1 U3928 ( .A0(N156), .A1(n3967), .B0(n3988), .B1(mem_wdata[18]), .Y(
        n2950) );
  AO22X1 U3929 ( .A0(N155), .A1(n3967), .B0(n3988), .B1(mem_wdata[19]), .Y(
        n2949) );
  AO22X1 U3930 ( .A0(N154), .A1(n3966), .B0(n3988), .B1(mem_wdata[20]), .Y(
        n2948) );
  AO22X1 U3931 ( .A0(N153), .A1(n3966), .B0(n3987), .B1(mem_wdata[21]), .Y(
        n2947) );
  AO22X1 U3932 ( .A0(N152), .A1(n3966), .B0(n3987), .B1(mem_wdata[22]), .Y(
        n2946) );
  AO22X1 U3933 ( .A0(N151), .A1(n3966), .B0(n3987), .B1(mem_wdata[23]), .Y(
        n2945) );
  AO22X1 U3934 ( .A0(N150), .A1(n3966), .B0(n3987), .B1(mem_wdata[24]), .Y(
        n2944) );
  AO22X1 U3935 ( .A0(N149), .A1(n3966), .B0(n3987), .B1(mem_wdata[25]), .Y(
        n2943) );
  AO22X1 U3936 ( .A0(N148), .A1(n3966), .B0(n3987), .B1(mem_wdata[26]), .Y(
        n2942) );
  AO22X1 U3937 ( .A0(N147), .A1(n3966), .B0(n3986), .B1(mem_wdata[27]), .Y(
        n2941) );
  AO22X1 U3938 ( .A0(N146), .A1(n3966), .B0(n3986), .B1(mem_wdata[28]), .Y(
        n2940) );
  AO22X1 U3939 ( .A0(N145), .A1(n3966), .B0(n3986), .B1(mem_wdata[29]), .Y(
        n2939) );
  AO22X1 U3940 ( .A0(N144), .A1(n3966), .B0(n3986), .B1(mem_wdata[30]), .Y(
        n2938) );
  AO22X1 U3941 ( .A0(N143), .A1(n3966), .B0(n3986), .B1(mem_wdata[31]), .Y(
        n2937) );
  AO22X1 U3942 ( .A0(N142), .A1(n3965), .B0(n3986), .B1(mem_wdata[32]), .Y(
        n2936) );
  AO22X1 U3943 ( .A0(N141), .A1(n3965), .B0(n3985), .B1(mem_wdata[33]), .Y(
        n2935) );
  AO22X1 U3944 ( .A0(N140), .A1(n3965), .B0(n3985), .B1(mem_wdata[34]), .Y(
        n2934) );
  AO22X1 U3945 ( .A0(N139), .A1(n3965), .B0(n3985), .B1(mem_wdata[35]), .Y(
        n2933) );
  AO22X1 U3946 ( .A0(N138), .A1(n3965), .B0(n3985), .B1(mem_wdata[36]), .Y(
        n2932) );
  AO22X1 U3947 ( .A0(N137), .A1(n3965), .B0(n3985), .B1(mem_wdata[37]), .Y(
        n2931) );
  AO22X1 U3948 ( .A0(N136), .A1(n3965), .B0(n3985), .B1(mem_wdata[38]), .Y(
        n2930) );
  AO22X1 U3949 ( .A0(N135), .A1(n3965), .B0(n3984), .B1(mem_wdata[39]), .Y(
        n2929) );
  AO22X1 U3950 ( .A0(N134), .A1(n3965), .B0(n3984), .B1(mem_wdata[40]), .Y(
        n2928) );
  AO22X1 U3951 ( .A0(N133), .A1(n3965), .B0(n3984), .B1(mem_wdata[41]), .Y(
        n2927) );
  AO22X1 U3952 ( .A0(N132), .A1(n3965), .B0(n3984), .B1(mem_wdata[42]), .Y(
        n2926) );
  AO22X1 U3953 ( .A0(N131), .A1(n3965), .B0(n3984), .B1(mem_wdata[43]), .Y(
        n2925) );
  AO22X1 U3954 ( .A0(N130), .A1(n3964), .B0(n3984), .B1(mem_wdata[44]), .Y(
        n2924) );
  AO22X1 U3955 ( .A0(N129), .A1(n3964), .B0(n3983), .B1(mem_wdata[45]), .Y(
        n2923) );
  AO22X1 U3956 ( .A0(N128), .A1(n3964), .B0(n3983), .B1(mem_wdata[46]), .Y(
        n2922) );
  AO22X1 U3957 ( .A0(N127), .A1(n3964), .B0(n3983), .B1(mem_wdata[47]), .Y(
        n2921) );
  AO22X1 U3958 ( .A0(N126), .A1(n3964), .B0(n3983), .B1(mem_wdata[48]), .Y(
        n2920) );
  AO22X1 U3959 ( .A0(N125), .A1(n3964), .B0(n3983), .B1(mem_wdata[49]), .Y(
        n2919) );
  AO22X1 U3960 ( .A0(N124), .A1(n3964), .B0(n3983), .B1(mem_wdata[50]), .Y(
        n2918) );
  AO22X1 U3961 ( .A0(N123), .A1(n3964), .B0(n3982), .B1(mem_wdata[51]), .Y(
        n2917) );
  AO22X1 U3962 ( .A0(N122), .A1(n3964), .B0(n3982), .B1(mem_wdata[52]), .Y(
        n2916) );
  AO22X1 U3963 ( .A0(N121), .A1(n3964), .B0(n3982), .B1(mem_wdata[53]), .Y(
        n2915) );
  AO22X1 U3964 ( .A0(N120), .A1(n3964), .B0(n3982), .B1(mem_wdata[54]), .Y(
        n2914) );
  AO22X1 U3965 ( .A0(N119), .A1(n3964), .B0(n3982), .B1(mem_wdata[55]), .Y(
        n2913) );
  AO22X1 U3966 ( .A0(N118), .A1(n3963), .B0(n3982), .B1(mem_wdata[56]), .Y(
        n2912) );
  AO22X1 U3967 ( .A0(N117), .A1(n3963), .B0(n3981), .B1(mem_wdata[57]), .Y(
        n2911) );
  AO22X1 U3968 ( .A0(N116), .A1(n3963), .B0(n3981), .B1(mem_wdata[58]), .Y(
        n2910) );
  AO22X1 U3969 ( .A0(N115), .A1(n3963), .B0(n3981), .B1(mem_wdata[59]), .Y(
        n2909) );
  AO22X1 U3970 ( .A0(N114), .A1(n3963), .B0(n3981), .B1(mem_wdata[60]), .Y(
        n2908) );
  AO22X1 U3971 ( .A0(N113), .A1(n3963), .B0(n3981), .B1(mem_wdata[61]), .Y(
        n2907) );
  AO22X1 U3972 ( .A0(N112), .A1(n3963), .B0(n3981), .B1(mem_wdata[62]), .Y(
        n2906) );
  AO22X1 U3973 ( .A0(N111), .A1(n3963), .B0(n3980), .B1(mem_wdata[63]), .Y(
        n2905) );
  AO22X1 U3974 ( .A0(N110), .A1(n3963), .B0(n3980), .B1(mem_wdata[64]), .Y(
        n2904) );
  AO22X1 U3975 ( .A0(N109), .A1(n3963), .B0(n3980), .B1(mem_wdata[65]), .Y(
        n2903) );
  AO22X1 U3976 ( .A0(N108), .A1(n3963), .B0(n3980), .B1(mem_wdata[66]), .Y(
        n2902) );
  AO22X1 U3977 ( .A0(N107), .A1(n3963), .B0(n3980), .B1(mem_wdata[67]), .Y(
        n2901) );
  AO22X1 U3978 ( .A0(N106), .A1(n3962), .B0(n3980), .B1(mem_wdata[68]), .Y(
        n2900) );
  AO22X1 U3979 ( .A0(N105), .A1(n3962), .B0(n3979), .B1(mem_wdata[69]), .Y(
        n2899) );
  AO22X1 U3980 ( .A0(N104), .A1(n3962), .B0(n3979), .B1(mem_wdata[70]), .Y(
        n2898) );
  AO22X1 U3981 ( .A0(N103), .A1(n3962), .B0(n3979), .B1(mem_wdata[71]), .Y(
        n2897) );
  AO22X1 U3982 ( .A0(N102), .A1(n3962), .B0(n3979), .B1(mem_wdata[72]), .Y(
        n2896) );
  AO22X1 U3983 ( .A0(N101), .A1(n3962), .B0(n3979), .B1(mem_wdata[73]), .Y(
        n2895) );
  AO22X1 U3984 ( .A0(N100), .A1(n3962), .B0(n3979), .B1(mem_wdata[74]), .Y(
        n2894) );
  AO22X1 U3985 ( .A0(N99), .A1(n3962), .B0(n3978), .B1(mem_wdata[75]), .Y(
        n2893) );
  AO22X1 U3986 ( .A0(N98), .A1(n3962), .B0(n3978), .B1(mem_wdata[76]), .Y(
        n2892) );
  AO22X1 U3987 ( .A0(N97), .A1(n3962), .B0(n3978), .B1(mem_wdata[77]), .Y(
        n2891) );
  AO22X1 U3988 ( .A0(N96), .A1(n3962), .B0(n3978), .B1(mem_wdata[78]), .Y(
        n2890) );
  AO22X1 U3989 ( .A0(N95), .A1(n3962), .B0(n3978), .B1(mem_wdata[79]), .Y(
        n2889) );
  AO22X1 U3990 ( .A0(N94), .A1(n3962), .B0(n3978), .B1(mem_wdata[80]), .Y(
        n2888) );
  AO22X1 U3991 ( .A0(N93), .A1(n3962), .B0(n3977), .B1(mem_wdata[81]), .Y(
        n2887) );
  AO22X1 U3992 ( .A0(N92), .A1(n3962), .B0(n3977), .B1(mem_wdata[82]), .Y(
        n2886) );
  AO22X1 U3993 ( .A0(N91), .A1(n3962), .B0(n3977), .B1(mem_wdata[83]), .Y(
        n2885) );
  AO22X1 U3994 ( .A0(N90), .A1(n3962), .B0(n3977), .B1(mem_wdata[84]), .Y(
        n2884) );
  AO22X1 U3995 ( .A0(N89), .A1(n3962), .B0(n3977), .B1(mem_wdata[85]), .Y(
        n2883) );
  AO22X1 U3996 ( .A0(N88), .A1(n3962), .B0(n3977), .B1(mem_wdata[86]), .Y(
        n2882) );
  AO22X1 U3997 ( .A0(N87), .A1(n3962), .B0(n3976), .B1(mem_wdata[87]), .Y(
        n2881) );
  AO22X1 U3998 ( .A0(N86), .A1(n3962), .B0(n3976), .B1(mem_wdata[88]), .Y(
        n2880) );
  AO22X1 U3999 ( .A0(N85), .A1(n3962), .B0(n3976), .B1(mem_wdata[89]), .Y(
        n2879) );
  AO22X1 U4000 ( .A0(N84), .A1(n3961), .B0(n3976), .B1(mem_wdata[90]), .Y(
        n2878) );
  AO22X1 U4001 ( .A0(N83), .A1(n3961), .B0(n3976), .B1(mem_wdata[91]), .Y(
        n2877) );
  AO22X1 U4002 ( .A0(N82), .A1(n3961), .B0(n3976), .B1(mem_wdata[92]), .Y(
        n2876) );
  AO22X1 U4003 ( .A0(N81), .A1(n3961), .B0(n3975), .B1(mem_wdata[93]), .Y(
        n2875) );
  AO22X1 U4004 ( .A0(N80), .A1(n3963), .B0(n3975), .B1(mem_wdata[94]), .Y(
        n2874) );
  AO22X1 U4005 ( .A0(N79), .A1(n3961), .B0(n3975), .B1(mem_wdata[95]), .Y(
        n2873) );
  AO22X1 U4006 ( .A0(N78), .A1(n3967), .B0(n3975), .B1(mem_wdata[96]), .Y(
        n2872) );
  AO22X1 U4007 ( .A0(N77), .A1(n3961), .B0(n3975), .B1(mem_wdata[97]), .Y(
        n2871) );
  AO22X1 U4008 ( .A0(N76), .A1(n3963), .B0(n3975), .B1(mem_wdata[98]), .Y(
        n2870) );
  AO22X1 U4009 ( .A0(N75), .A1(n3965), .B0(n3974), .B1(mem_wdata[99]), .Y(
        n2869) );
  AO22X1 U4010 ( .A0(N74), .A1(n3961), .B0(n3974), .B1(mem_wdata[100]), .Y(
        n2868) );
  AO22X1 U4011 ( .A0(N73), .A1(n3963), .B0(n3974), .B1(mem_wdata[101]), .Y(
        n2867) );
  AO22X1 U4012 ( .A0(N72), .A1(n3966), .B0(n3974), .B1(mem_wdata[102]), .Y(
        n2866) );
  AO22X1 U4013 ( .A0(N71), .A1(n3966), .B0(n3974), .B1(mem_wdata[103]), .Y(
        n2865) );
  AO22X1 U4014 ( .A0(N70), .A1(n3963), .B0(n3974), .B1(mem_wdata[104]), .Y(
        n2864) );
  AO22X1 U4015 ( .A0(N69), .A1(n3967), .B0(n3973), .B1(mem_wdata[105]), .Y(
        n2863) );
  AO22X1 U4016 ( .A0(N68), .A1(n3965), .B0(n3973), .B1(mem_wdata[106]), .Y(
        n2862) );
  AO22X1 U4017 ( .A0(N67), .A1(n3966), .B0(n3973), .B1(mem_wdata[107]), .Y(
        n2861) );
  AO22X1 U4018 ( .A0(N66), .A1(n3968), .B0(n3973), .B1(mem_wdata[108]), .Y(
        n2860) );
  AO22X1 U4019 ( .A0(N65), .A1(n3961), .B0(n3973), .B1(mem_wdata[109]), .Y(
        n2859) );
  AO22X1 U4020 ( .A0(N64), .A1(n3963), .B0(n3973), .B1(mem_wdata[110]), .Y(
        n2858) );
  AO22X1 U4021 ( .A0(N63), .A1(n3967), .B0(n3972), .B1(mem_wdata[111]), .Y(
        n2857) );
  AO22X1 U4022 ( .A0(N62), .A1(n3965), .B0(n3972), .B1(mem_wdata[112]), .Y(
        n2856) );
  AO22X1 U4023 ( .A0(N61), .A1(n3966), .B0(n3972), .B1(mem_wdata[113]), .Y(
        n2855) );
  AO22X1 U4024 ( .A0(N60), .A1(n3968), .B0(n3972), .B1(mem_wdata[114]), .Y(
        n2854) );
  AO22X1 U4025 ( .A0(N59), .A1(n3961), .B0(n3972), .B1(mem_wdata[115]), .Y(
        n2853) );
  AO22X1 U4026 ( .A0(N58), .A1(n3961), .B0(n3972), .B1(mem_wdata[116]), .Y(
        n2852) );
  AO22X1 U4027 ( .A0(N57), .A1(n3961), .B0(n3997), .B1(mem_wdata[117]), .Y(
        n2851) );
  AO22X1 U4028 ( .A0(N56), .A1(n3961), .B0(n3997), .B1(mem_wdata[118]), .Y(
        n2850) );
  AO22X1 U4029 ( .A0(N55), .A1(n3961), .B0(n3997), .B1(mem_wdata[119]), .Y(
        n2849) );
  AO22X1 U4030 ( .A0(N54), .A1(n3961), .B0(n3997), .B1(mem_wdata[120]), .Y(
        n2848) );
  AO22X1 U4031 ( .A0(N53), .A1(n3961), .B0(n3997), .B1(mem_wdata[121]), .Y(
        n2847) );
  AO22X1 U4032 ( .A0(N52), .A1(n3961), .B0(n3971), .B1(mem_wdata[122]), .Y(
        n2846) );
  AO22X1 U4033 ( .A0(N51), .A1(n3961), .B0(n3991), .B1(mem_wdata[123]), .Y(
        n2845) );
  AO22X1 U4034 ( .A0(N50), .A1(n3961), .B0(n3970), .B1(mem_wdata[124]), .Y(
        n2844) );
  AO22X1 U4035 ( .A0(N49), .A1(n3961), .B0(n3970), .B1(mem_wdata[125]), .Y(
        n2843) );
  AO22X1 U4036 ( .A0(N48), .A1(n3961), .B0(n3969), .B1(mem_wdata[126]), .Y(
        n2842) );
  AO22X1 U4037 ( .A0(N47), .A1(n3961), .B0(n3991), .B1(mem_wdata[127]), .Y(
        n2841) );
  OA22X1 U4038 ( .A0(rw_status), .A1(n198), .B0(n199), .B1(n200), .Y(n3282) );
  CLKINVX1 U4039 ( .A(n3282), .Y(n197) );
  MXI2X1 U4040 ( .A(n3466), .B(n3467), .S0(n3665), .Y(N110) );
  MXI4X1 U4041 ( .A(\block[0][2][0] ), .B(\block[1][2][0] ), .C(
        \block[2][2][0] ), .D(\block[3][2][0] ), .S0(n3616), .S1(n3645), .Y(
        n3466) );
  MXI4X1 U4042 ( .A(\block[4][2][0] ), .B(\block[5][2][0] ), .C(
        \block[6][2][0] ), .D(\block[7][2][0] ), .S0(n3609), .S1(n3645), .Y(
        n3467) );
  MXI2X1 U4043 ( .A(n3464), .B(n3465), .S0(n3662), .Y(N109) );
  MXI4X1 U4044 ( .A(\block[0][2][1] ), .B(\block[1][2][1] ), .C(
        \block[2][2][1] ), .D(\block[3][2][1] ), .S0(n3615), .S1(n3645), .Y(
        n3464) );
  MXI4X1 U4045 ( .A(\block[4][2][1] ), .B(\block[5][2][1] ), .C(
        \block[6][2][1] ), .D(\block[7][2][1] ), .S0(n3615), .S1(n3645), .Y(
        n3465) );
  MXI2X1 U4046 ( .A(n3462), .B(n3463), .S0(n3661), .Y(N108) );
  MXI4X1 U4047 ( .A(\block[0][2][2] ), .B(\block[1][2][2] ), .C(
        \block[2][2][2] ), .D(\block[3][2][2] ), .S0(n3615), .S1(n3644), .Y(
        n3462) );
  MXI4X1 U4048 ( .A(\block[4][2][2] ), .B(\block[5][2][2] ), .C(
        \block[6][2][2] ), .D(\block[7][2][2] ), .S0(n3615), .S1(n3644), .Y(
        n3463) );
  MXI2X1 U4049 ( .A(n3460), .B(n3461), .S0(n3660), .Y(N107) );
  MXI4X1 U4050 ( .A(\block[0][2][3] ), .B(\block[1][2][3] ), .C(
        \block[2][2][3] ), .D(\block[3][2][3] ), .S0(n3615), .S1(n3644), .Y(
        n3460) );
  MXI4X1 U4051 ( .A(\block[4][2][3] ), .B(\block[5][2][3] ), .C(
        \block[6][2][3] ), .D(\block[7][2][3] ), .S0(n3615), .S1(n3644), .Y(
        n3461) );
  MXI2X1 U4052 ( .A(n3458), .B(n3459), .S0(n3662), .Y(N106) );
  MXI4X1 U4053 ( .A(\block[0][2][4] ), .B(\block[1][2][4] ), .C(
        \block[2][2][4] ), .D(\block[3][2][4] ), .S0(n3615), .S1(n3644), .Y(
        n3458) );
  MXI4X1 U4054 ( .A(\block[4][2][4] ), .B(\block[5][2][4] ), .C(
        \block[6][2][4] ), .D(\block[7][2][4] ), .S0(n3615), .S1(n3644), .Y(
        n3459) );
  MXI2X1 U4055 ( .A(n3456), .B(n3457), .S0(n3661), .Y(N105) );
  MXI4X1 U4056 ( .A(\block[0][2][5] ), .B(\block[1][2][5] ), .C(
        \block[2][2][5] ), .D(\block[3][2][5] ), .S0(n3615), .S1(n3644), .Y(
        n3456) );
  MXI4X1 U4057 ( .A(\block[4][2][5] ), .B(\block[5][2][5] ), .C(
        \block[6][2][5] ), .D(\block[7][2][5] ), .S0(n3615), .S1(n3644), .Y(
        n3457) );
  MXI2X1 U4058 ( .A(n3454), .B(n3455), .S0(n3660), .Y(N104) );
  MXI4X1 U4059 ( .A(\block[0][2][6] ), .B(\block[1][2][6] ), .C(
        \block[2][2][6] ), .D(\block[3][2][6] ), .S0(n3615), .S1(n3644), .Y(
        n3454) );
  MXI4X1 U4060 ( .A(\block[4][2][6] ), .B(\block[5][2][6] ), .C(
        \block[6][2][6] ), .D(\block[7][2][6] ), .S0(n3615), .S1(n3644), .Y(
        n3455) );
  MXI2X1 U4061 ( .A(n3452), .B(n3453), .S0(n3666), .Y(N103) );
  MXI4X1 U4062 ( .A(\block[0][2][7] ), .B(\block[1][2][7] ), .C(
        \block[2][2][7] ), .D(\block[3][2][7] ), .S0(n3615), .S1(n3644), .Y(
        n3452) );
  MXI4X1 U4063 ( .A(\block[4][2][7] ), .B(\block[5][2][7] ), .C(
        \block[6][2][7] ), .D(\block[7][2][7] ), .S0(n3614), .S1(n3644), .Y(
        n3453) );
  MXI2X1 U4064 ( .A(n3450), .B(n3451), .S0(n3662), .Y(N102) );
  MXI4X1 U4065 ( .A(\block[0][2][8] ), .B(\block[1][2][8] ), .C(
        \block[2][2][8] ), .D(\block[3][2][8] ), .S0(n3614), .S1(n3643), .Y(
        n3450) );
  MXI4X1 U4066 ( .A(\block[4][2][8] ), .B(\block[5][2][8] ), .C(
        \block[6][2][8] ), .D(\block[7][2][8] ), .S0(n3614), .S1(n3643), .Y(
        n3451) );
  MXI2X1 U4067 ( .A(n3448), .B(n3449), .S0(n3662), .Y(N101) );
  MXI4X1 U4068 ( .A(\block[0][2][9] ), .B(\block[1][2][9] ), .C(
        \block[2][2][9] ), .D(\block[3][2][9] ), .S0(n3614), .S1(n3643), .Y(
        n3448) );
  MXI4X1 U4069 ( .A(\block[4][2][9] ), .B(\block[5][2][9] ), .C(
        \block[6][2][9] ), .D(\block[7][2][9] ), .S0(n3614), .S1(n3643), .Y(
        n3449) );
  MXI2X1 U4070 ( .A(n3446), .B(n3447), .S0(n3662), .Y(N100) );
  MXI4X1 U4071 ( .A(\block[0][2][10] ), .B(\block[1][2][10] ), .C(
        \block[2][2][10] ), .D(\block[3][2][10] ), .S0(n3614), .S1(n3643), .Y(
        n3446) );
  MXI4X1 U4072 ( .A(\block[4][2][10] ), .B(\block[5][2][10] ), .C(
        \block[6][2][10] ), .D(\block[7][2][10] ), .S0(n3614), .S1(n3643), .Y(
        n3447) );
  MXI2X1 U4073 ( .A(n3444), .B(n3445), .S0(n3662), .Y(N99) );
  MXI4X1 U4074 ( .A(\block[0][2][11] ), .B(\block[1][2][11] ), .C(
        \block[2][2][11] ), .D(\block[3][2][11] ), .S0(n3614), .S1(n3643), .Y(
        n3444) );
  MXI4X1 U4075 ( .A(\block[4][2][11] ), .B(\block[5][2][11] ), .C(
        \block[6][2][11] ), .D(\block[7][2][11] ), .S0(n3614), .S1(n3643), .Y(
        n3445) );
  MXI2X1 U4076 ( .A(n3442), .B(n3443), .S0(n3662), .Y(N98) );
  MXI4X1 U4077 ( .A(\block[0][2][12] ), .B(\block[1][2][12] ), .C(
        \block[2][2][12] ), .D(\block[3][2][12] ), .S0(n3614), .S1(n3643), .Y(
        n3442) );
  MXI4X1 U4078 ( .A(\block[4][2][12] ), .B(\block[5][2][12] ), .C(
        \block[6][2][12] ), .D(\block[7][2][12] ), .S0(n3614), .S1(n3643), .Y(
        n3443) );
  MXI2X1 U4079 ( .A(n3440), .B(n3441), .S0(n3662), .Y(N97) );
  MXI4X1 U4080 ( .A(\block[0][2][13] ), .B(\block[1][2][13] ), .C(
        \block[2][2][13] ), .D(\block[3][2][13] ), .S0(n3614), .S1(n3643), .Y(
        n3440) );
  MXI4X1 U4081 ( .A(\block[4][2][13] ), .B(\block[5][2][13] ), .C(
        \block[6][2][13] ), .D(\block[7][2][13] ), .S0(n3614), .S1(n3643), .Y(
        n3441) );
  MXI2X1 U4082 ( .A(n3438), .B(n3439), .S0(n3662), .Y(N96) );
  MXI4X1 U4083 ( .A(\block[0][2][14] ), .B(\block[1][2][14] ), .C(
        \block[2][2][14] ), .D(\block[3][2][14] ), .S0(n3613), .S1(n3642), .Y(
        n3438) );
  MXI4X1 U4084 ( .A(\block[4][2][14] ), .B(\block[5][2][14] ), .C(
        \block[6][2][14] ), .D(\block[7][2][14] ), .S0(n3613), .S1(n3642), .Y(
        n3439) );
  MXI2X1 U4085 ( .A(n3436), .B(n3437), .S0(n3662), .Y(N95) );
  MXI4X1 U4086 ( .A(\block[0][2][15] ), .B(\block[1][2][15] ), .C(
        \block[2][2][15] ), .D(\block[3][2][15] ), .S0(n3613), .S1(n3642), .Y(
        n3436) );
  MXI4X1 U4087 ( .A(\block[4][2][15] ), .B(\block[5][2][15] ), .C(
        \block[6][2][15] ), .D(\block[7][2][15] ), .S0(n3613), .S1(n3642), .Y(
        n3437) );
  MXI2X1 U4088 ( .A(n3434), .B(n3435), .S0(n3662), .Y(N94) );
  MXI4X1 U4089 ( .A(\block[0][2][16] ), .B(\block[1][2][16] ), .C(
        \block[2][2][16] ), .D(\block[3][2][16] ), .S0(n3613), .S1(n3642), .Y(
        n3434) );
  MXI4X1 U4090 ( .A(\block[4][2][16] ), .B(\block[5][2][16] ), .C(
        \block[6][2][16] ), .D(\block[7][2][16] ), .S0(n3613), .S1(n3642), .Y(
        n3435) );
  MXI2X1 U4091 ( .A(n3432), .B(n3433), .S0(n3662), .Y(N93) );
  MXI4X1 U4092 ( .A(\block[0][2][17] ), .B(\block[1][2][17] ), .C(
        \block[2][2][17] ), .D(\block[3][2][17] ), .S0(n3613), .S1(n3642), .Y(
        n3432) );
  MXI4X1 U4093 ( .A(\block[4][2][17] ), .B(\block[5][2][17] ), .C(
        \block[6][2][17] ), .D(\block[7][2][17] ), .S0(n3613), .S1(n3642), .Y(
        n3433) );
  MXI2X1 U4094 ( .A(n3430), .B(n3431), .S0(n3662), .Y(N92) );
  MXI4X1 U4095 ( .A(\block[0][2][18] ), .B(\block[1][2][18] ), .C(
        \block[2][2][18] ), .D(\block[3][2][18] ), .S0(n3613), .S1(n3642), .Y(
        n3430) );
  MXI4X1 U4096 ( .A(\block[4][2][18] ), .B(\block[5][2][18] ), .C(
        \block[6][2][18] ), .D(\block[7][2][18] ), .S0(n3613), .S1(n3642), .Y(
        n3431) );
  MXI2X1 U4097 ( .A(n3428), .B(n3429), .S0(n3662), .Y(N91) );
  MXI4X1 U4098 ( .A(\block[0][2][19] ), .B(\block[1][2][19] ), .C(
        \block[2][2][19] ), .D(\block[3][2][19] ), .S0(n3613), .S1(n3642), .Y(
        n3428) );
  MXI4X1 U4099 ( .A(\block[4][2][19] ), .B(\block[5][2][19] ), .C(
        \block[6][2][19] ), .D(\block[7][2][19] ), .S0(n3613), .S1(n3642), .Y(
        n3429) );
  MXI2X1 U4100 ( .A(n3426), .B(n3427), .S0(n3661), .Y(N90) );
  MXI4X1 U4101 ( .A(\block[0][2][20] ), .B(\block[1][2][20] ), .C(
        \block[2][2][20] ), .D(\block[3][2][20] ), .S0(n3613), .S1(n3641), .Y(
        n3426) );
  MXI4X1 U4102 ( .A(\block[4][2][20] ), .B(\block[5][2][20] ), .C(
        \block[6][2][20] ), .D(\block[7][2][20] ), .S0(n3612), .S1(n3641), .Y(
        n3427) );
  MXI2X1 U4103 ( .A(n3424), .B(n3425), .S0(n3661), .Y(N89) );
  MXI4X1 U4104 ( .A(\block[0][2][21] ), .B(\block[1][2][21] ), .C(
        \block[2][2][21] ), .D(\block[3][2][21] ), .S0(n3612), .S1(n3641), .Y(
        n3424) );
  MXI4X1 U4105 ( .A(\block[4][2][21] ), .B(\block[5][2][21] ), .C(
        \block[6][2][21] ), .D(\block[7][2][21] ), .S0(n3612), .S1(n3641), .Y(
        n3425) );
  MXI2X1 U4106 ( .A(n3422), .B(n3423), .S0(n3661), .Y(N88) );
  MXI4X1 U4107 ( .A(\block[0][2][22] ), .B(\block[1][2][22] ), .C(
        \block[2][2][22] ), .D(\block[3][2][22] ), .S0(n3612), .S1(n3641), .Y(
        n3422) );
  MXI4X1 U4108 ( .A(\block[4][2][22] ), .B(\block[5][2][22] ), .C(
        \block[6][2][22] ), .D(\block[7][2][22] ), .S0(n3612), .S1(n3641), .Y(
        n3423) );
  MXI2X1 U4109 ( .A(n3420), .B(n3421), .S0(n3661), .Y(N87) );
  MXI4X1 U4110 ( .A(\block[0][2][23] ), .B(\block[1][2][23] ), .C(
        \block[2][2][23] ), .D(\block[3][2][23] ), .S0(n3612), .S1(n3641), .Y(
        n3420) );
  MXI4X1 U4111 ( .A(\block[4][2][23] ), .B(\block[5][2][23] ), .C(
        \block[6][2][23] ), .D(\block[7][2][23] ), .S0(n3612), .S1(n3641), .Y(
        n3421) );
  MXI2X1 U4112 ( .A(n3418), .B(n3419), .S0(n3661), .Y(N86) );
  MXI4X1 U4113 ( .A(\block[0][2][24] ), .B(\block[1][2][24] ), .C(
        \block[2][2][24] ), .D(\block[3][2][24] ), .S0(n3612), .S1(n3641), .Y(
        n3418) );
  MXI4X1 U4114 ( .A(\block[4][2][24] ), .B(\block[5][2][24] ), .C(
        \block[6][2][24] ), .D(\block[7][2][24] ), .S0(n3612), .S1(n3641), .Y(
        n3419) );
  MXI2X1 U4115 ( .A(n3416), .B(n3417), .S0(n3661), .Y(N85) );
  MXI4X1 U4116 ( .A(\block[0][2][25] ), .B(\block[1][2][25] ), .C(
        \block[2][2][25] ), .D(\block[3][2][25] ), .S0(n3612), .S1(n3641), .Y(
        n3416) );
  MXI4X1 U4117 ( .A(\block[4][2][25] ), .B(\block[5][2][25] ), .C(
        \block[6][2][25] ), .D(\block[7][2][25] ), .S0(n3612), .S1(n3641), .Y(
        n3417) );
  MXI2X1 U4118 ( .A(n3414), .B(n3415), .S0(n3661), .Y(N84) );
  MXI4X1 U4119 ( .A(\block[0][2][26] ), .B(\block[1][2][26] ), .C(
        \block[2][2][26] ), .D(\block[3][2][26] ), .S0(n3612), .S1(n3640), .Y(
        n3414) );
  MXI4X1 U4120 ( .A(\block[4][2][26] ), .B(\block[5][2][26] ), .C(
        \block[6][2][26] ), .D(\block[7][2][26] ), .S0(n3612), .S1(n3640), .Y(
        n3415) );
  MXI2X1 U4121 ( .A(n3412), .B(n3413), .S0(n3661), .Y(N83) );
  MXI4X1 U4122 ( .A(\block[0][2][27] ), .B(\block[1][2][27] ), .C(
        \block[2][2][27] ), .D(\block[3][2][27] ), .S0(n3611), .S1(n3640), .Y(
        n3412) );
  MXI4X1 U4123 ( .A(\block[4][2][27] ), .B(\block[5][2][27] ), .C(
        \block[6][2][27] ), .D(\block[7][2][27] ), .S0(n3611), .S1(n3640), .Y(
        n3413) );
  MXI2X1 U4124 ( .A(n3410), .B(n3411), .S0(n3661), .Y(N82) );
  MXI4X1 U4125 ( .A(\block[0][2][28] ), .B(\block[1][2][28] ), .C(
        \block[2][2][28] ), .D(\block[3][2][28] ), .S0(n3611), .S1(n3640), .Y(
        n3410) );
  MXI4X1 U4126 ( .A(\block[4][2][28] ), .B(\block[5][2][28] ), .C(
        \block[6][2][28] ), .D(\block[7][2][28] ), .S0(n3611), .S1(n3640), .Y(
        n3411) );
  MXI2X1 U4127 ( .A(n3408), .B(n3409), .S0(n3661), .Y(N81) );
  MXI4X1 U4128 ( .A(\block[0][2][29] ), .B(\block[1][2][29] ), .C(
        \block[2][2][29] ), .D(\block[3][2][29] ), .S0(n3611), .S1(n3640), .Y(
        n3408) );
  MXI4X1 U4129 ( .A(\block[4][2][29] ), .B(\block[5][2][29] ), .C(
        \block[6][2][29] ), .D(\block[7][2][29] ), .S0(n3611), .S1(n3640), .Y(
        n3409) );
  MXI2X1 U4130 ( .A(n3406), .B(n3407), .S0(n3661), .Y(N80) );
  MXI4X1 U4131 ( .A(\block[0][2][30] ), .B(\block[1][2][30] ), .C(
        \block[2][2][30] ), .D(\block[3][2][30] ), .S0(n3611), .S1(n3640), .Y(
        n3406) );
  MXI4X1 U4132 ( .A(\block[4][2][30] ), .B(\block[5][2][30] ), .C(
        \block[6][2][30] ), .D(\block[7][2][30] ), .S0(n3611), .S1(n3640), .Y(
        n3407) );
  MXI2X1 U4133 ( .A(n3404), .B(n3405), .S0(n3661), .Y(N79) );
  MXI4X1 U4134 ( .A(\block[0][2][31] ), .B(\block[1][2][31] ), .C(
        \block[2][2][31] ), .D(\block[3][2][31] ), .S0(n3611), .S1(n3640), .Y(
        n3404) );
  MXI4X1 U4135 ( .A(\block[4][2][31] ), .B(\block[5][2][31] ), .C(
        \block[6][2][31] ), .D(\block[7][2][31] ), .S0(n3611), .S1(n3640), .Y(
        n3405) );
  MXI2X1 U4136 ( .A(n3594), .B(n3595), .S0(n3666), .Y(N174) );
  MXI4X1 U4137 ( .A(\block[0][0][0] ), .B(\block[1][0][0] ), .C(
        \block[2][0][0] ), .D(\block[3][0][0] ), .S0(n3622), .S1(n3654), .Y(
        n3594) );
  MXI4X1 U4138 ( .A(\block[4][0][0] ), .B(\block[5][0][0] ), .C(
        \block[6][0][0] ), .D(\block[7][0][0] ), .S0(n3622), .S1(n3654), .Y(
        n3595) );
  MXI2X1 U4139 ( .A(n3592), .B(n3593), .S0(n3666), .Y(N173) );
  MXI4X1 U4140 ( .A(\block[0][0][1] ), .B(\block[1][0][1] ), .C(
        \block[2][0][1] ), .D(\block[3][0][1] ), .S0(n3622), .S1(n3654), .Y(
        n3592) );
  MXI4X1 U4141 ( .A(\block[4][0][1] ), .B(\block[5][0][1] ), .C(
        \block[6][0][1] ), .D(\block[7][0][1] ), .S0(n3622), .S1(n3654), .Y(
        n3593) );
  MXI2X1 U4142 ( .A(n3590), .B(n3591), .S0(n3666), .Y(N172) );
  MXI4X1 U4143 ( .A(\block[0][0][2] ), .B(\block[1][0][2] ), .C(
        \block[2][0][2] ), .D(\block[3][0][2] ), .S0(n3622), .S1(n3654), .Y(
        n3590) );
  MXI4X1 U4144 ( .A(\block[4][0][2] ), .B(\block[5][0][2] ), .C(
        \block[6][0][2] ), .D(\block[7][0][2] ), .S0(n3622), .S1(n3654), .Y(
        n3591) );
  MXI2X1 U4145 ( .A(n3588), .B(n3589), .S0(n3666), .Y(N171) );
  MXI4X1 U4146 ( .A(\block[0][0][3] ), .B(\block[1][0][3] ), .C(
        \block[2][0][3] ), .D(\block[3][0][3] ), .S0(n3622), .S1(n3654), .Y(
        n3588) );
  MXI4X1 U4147 ( .A(\block[4][0][3] ), .B(\block[5][0][3] ), .C(
        \block[6][0][3] ), .D(\block[7][0][3] ), .S0(n3622), .S1(n3654), .Y(
        n3589) );
  MXI2X1 U4148 ( .A(n3586), .B(n3587), .S0(n3666), .Y(N170) );
  MXI4X1 U4149 ( .A(\block[0][0][4] ), .B(\block[1][0][4] ), .C(
        \block[2][0][4] ), .D(\block[3][0][4] ), .S0(n3622), .S1(n3654), .Y(
        n3586) );
  MXI4X1 U4150 ( .A(\block[4][0][4] ), .B(\block[5][0][4] ), .C(
        \block[6][0][4] ), .D(\block[7][0][4] ), .S0(n3622), .S1(n3654), .Y(
        n3587) );
  MXI2X1 U4151 ( .A(n3584), .B(n3585), .S0(n3666), .Y(N169) );
  MXI4X1 U4152 ( .A(\block[0][0][5] ), .B(\block[1][0][5] ), .C(
        \block[2][0][5] ), .D(\block[3][0][5] ), .S0(n3622), .S1(n3654), .Y(
        n3584) );
  MXI4X1 U4153 ( .A(\block[4][0][5] ), .B(\block[5][0][5] ), .C(
        \block[6][0][5] ), .D(\block[7][0][5] ), .S0(n3622), .S1(n3654), .Y(
        n3585) );
  MXI2X1 U4154 ( .A(n3582), .B(n3583), .S0(n3666), .Y(N168) );
  MXI4X1 U4155 ( .A(\block[0][0][6] ), .B(\block[1][0][6] ), .C(
        \block[2][0][6] ), .D(\block[3][0][6] ), .S0(n3622), .S1(n3653), .Y(
        n3582) );
  MXI4X1 U4156 ( .A(\block[4][0][6] ), .B(\block[5][0][6] ), .C(
        \block[6][0][6] ), .D(\block[7][0][6] ), .S0(n3621), .S1(n3653), .Y(
        n3583) );
  MXI2X1 U4157 ( .A(n3580), .B(n3581), .S0(n3666), .Y(N167) );
  MXI4X1 U4158 ( .A(\block[0][0][7] ), .B(\block[1][0][7] ), .C(
        \block[2][0][7] ), .D(\block[3][0][7] ), .S0(n3621), .S1(n3653), .Y(
        n3580) );
  MXI4X1 U4159 ( .A(\block[4][0][7] ), .B(\block[5][0][7] ), .C(
        \block[6][0][7] ), .D(\block[7][0][7] ), .S0(n3621), .S1(n3653), .Y(
        n3581) );
  MXI2X1 U4160 ( .A(n3578), .B(n3579), .S0(n3666), .Y(N166) );
  MXI4X1 U4161 ( .A(\block[0][0][8] ), .B(\block[1][0][8] ), .C(
        \block[2][0][8] ), .D(\block[3][0][8] ), .S0(n3621), .S1(n3653), .Y(
        n3578) );
  MXI4X1 U4162 ( .A(\block[4][0][8] ), .B(\block[5][0][8] ), .C(
        \block[6][0][8] ), .D(\block[7][0][8] ), .S0(n3621), .S1(n3653), .Y(
        n3579) );
  MXI2X1 U4163 ( .A(n3576), .B(n3577), .S0(n3666), .Y(N165) );
  MXI4X1 U4164 ( .A(\block[0][0][9] ), .B(\block[1][0][9] ), .C(
        \block[2][0][9] ), .D(\block[3][0][9] ), .S0(n3621), .S1(n3653), .Y(
        n3576) );
  MXI4X1 U4165 ( .A(\block[4][0][9] ), .B(\block[5][0][9] ), .C(
        \block[6][0][9] ), .D(\block[7][0][9] ), .S0(n3621), .S1(n3653), .Y(
        n3577) );
  MXI2X1 U4166 ( .A(n3574), .B(n3575), .S0(n3666), .Y(N164) );
  MXI4X1 U4167 ( .A(\block[0][0][10] ), .B(\block[1][0][10] ), .C(
        \block[2][0][10] ), .D(\block[3][0][10] ), .S0(n3621), .S1(n3653), .Y(
        n3574) );
  MXI4X1 U4168 ( .A(\block[4][0][10] ), .B(\block[5][0][10] ), .C(
        \block[6][0][10] ), .D(\block[7][0][10] ), .S0(n3621), .S1(n3653), .Y(
        n3575) );
  MXI2X1 U4169 ( .A(n3572), .B(n3573), .S0(n3666), .Y(N163) );
  MXI4X1 U4170 ( .A(\block[0][0][11] ), .B(\block[1][0][11] ), .C(
        \block[2][0][11] ), .D(\block[3][0][11] ), .S0(n3621), .S1(n3653), .Y(
        n3572) );
  MXI4X1 U4171 ( .A(\block[4][0][11] ), .B(\block[5][0][11] ), .C(
        \block[6][0][11] ), .D(\block[7][0][11] ), .S0(n3621), .S1(n3653), .Y(
        n3573) );
  MXI2X1 U4172 ( .A(n3570), .B(n3571), .S0(n3665), .Y(N162) );
  MXI4X1 U4173 ( .A(\block[0][0][12] ), .B(\block[1][0][12] ), .C(
        \block[2][0][12] ), .D(\block[3][0][12] ), .S0(n3621), .S1(n3652), .Y(
        n3570) );
  MXI4X1 U4174 ( .A(\block[4][0][12] ), .B(\block[5][0][12] ), .C(
        \block[6][0][12] ), .D(\block[7][0][12] ), .S0(n3621), .S1(n3652), .Y(
        n3571) );
  MXI2X1 U4175 ( .A(n3568), .B(n3569), .S0(n3665), .Y(N161) );
  MXI4X1 U4176 ( .A(\block[0][0][13] ), .B(\block[1][0][13] ), .C(
        \block[2][0][13] ), .D(\block[3][0][13] ), .S0(n3620), .S1(n3652), .Y(
        n3568) );
  MXI4X1 U4177 ( .A(\block[4][0][13] ), .B(\block[5][0][13] ), .C(
        \block[6][0][13] ), .D(\block[7][0][13] ), .S0(n3620), .S1(n3652), .Y(
        n3569) );
  MXI2X1 U4178 ( .A(n3566), .B(n3567), .S0(n3665), .Y(N160) );
  MXI4X1 U4179 ( .A(\block[0][0][14] ), .B(\block[1][0][14] ), .C(
        \block[2][0][14] ), .D(\block[3][0][14] ), .S0(n3620), .S1(n3652), .Y(
        n3566) );
  MXI4X1 U4180 ( .A(\block[4][0][14] ), .B(\block[5][0][14] ), .C(
        \block[6][0][14] ), .D(\block[7][0][14] ), .S0(n3620), .S1(n3652), .Y(
        n3567) );
  MXI2X1 U4181 ( .A(n3564), .B(n3565), .S0(n3665), .Y(N159) );
  MXI4X1 U4182 ( .A(\block[0][0][15] ), .B(\block[1][0][15] ), .C(
        \block[2][0][15] ), .D(\block[3][0][15] ), .S0(n3620), .S1(n3652), .Y(
        n3564) );
  MXI4X1 U4183 ( .A(\block[4][0][15] ), .B(\block[5][0][15] ), .C(
        \block[6][0][15] ), .D(\block[7][0][15] ), .S0(n3620), .S1(n3652), .Y(
        n3565) );
  MXI2X1 U4184 ( .A(n3562), .B(n3563), .S0(n3665), .Y(N158) );
  MXI4X1 U4185 ( .A(\block[0][0][16] ), .B(\block[1][0][16] ), .C(
        \block[2][0][16] ), .D(\block[3][0][16] ), .S0(n3620), .S1(n3652), .Y(
        n3562) );
  MXI4X1 U4186 ( .A(\block[4][0][16] ), .B(\block[5][0][16] ), .C(
        \block[6][0][16] ), .D(\block[7][0][16] ), .S0(n3620), .S1(n3652), .Y(
        n3563) );
  MXI2X1 U4187 ( .A(n3560), .B(n3561), .S0(n3665), .Y(N157) );
  MXI4X1 U4188 ( .A(\block[0][0][17] ), .B(\block[1][0][17] ), .C(
        \block[2][0][17] ), .D(\block[3][0][17] ), .S0(n3620), .S1(n3652), .Y(
        n3560) );
  MXI4X1 U4189 ( .A(\block[4][0][17] ), .B(\block[5][0][17] ), .C(
        \block[6][0][17] ), .D(\block[7][0][17] ), .S0(n3620), .S1(n3652), .Y(
        n3561) );
  MXI2X1 U4190 ( .A(n3558), .B(n3559), .S0(n3665), .Y(N156) );
  MXI4X1 U4191 ( .A(\block[0][0][18] ), .B(\block[1][0][18] ), .C(
        \block[2][0][18] ), .D(\block[3][0][18] ), .S0(n3620), .S1(n3651), .Y(
        n3558) );
  MXI4X1 U4192 ( .A(\block[4][0][18] ), .B(\block[5][0][18] ), .C(
        \block[6][0][18] ), .D(\block[7][0][18] ), .S0(n3620), .S1(n3651), .Y(
        n3559) );
  MXI2X1 U4193 ( .A(n3556), .B(n3557), .S0(n3665), .Y(N155) );
  MXI4X1 U4194 ( .A(\block[0][0][19] ), .B(\block[1][0][19] ), .C(
        \block[2][0][19] ), .D(\block[3][0][19] ), .S0(n3620), .S1(n3651), .Y(
        n3556) );
  MXI4X1 U4195 ( .A(\block[4][0][19] ), .B(\block[5][0][19] ), .C(
        \block[6][0][19] ), .D(\block[7][0][19] ), .S0(n3619), .S1(n3651), .Y(
        n3557) );
  MXI2X1 U4196 ( .A(n3554), .B(n3555), .S0(n3665), .Y(N154) );
  MXI4X1 U4197 ( .A(\block[0][0][20] ), .B(\block[1][0][20] ), .C(
        \block[2][0][20] ), .D(\block[3][0][20] ), .S0(n3619), .S1(n3651), .Y(
        n3554) );
  MXI4X1 U4198 ( .A(\block[4][0][20] ), .B(\block[5][0][20] ), .C(
        \block[6][0][20] ), .D(\block[7][0][20] ), .S0(n3619), .S1(n3651), .Y(
        n3555) );
  MXI2X1 U4199 ( .A(n3552), .B(n3553), .S0(n3665), .Y(N153) );
  MXI4X1 U4200 ( .A(\block[0][0][21] ), .B(\block[1][0][21] ), .C(
        \block[2][0][21] ), .D(\block[3][0][21] ), .S0(n3619), .S1(n3651), .Y(
        n3552) );
  MXI4X1 U4201 ( .A(\block[4][0][21] ), .B(\block[5][0][21] ), .C(
        \block[6][0][21] ), .D(\block[7][0][21] ), .S0(n3619), .S1(n3651), .Y(
        n3553) );
  MXI2X1 U4202 ( .A(n3550), .B(n3551), .S0(n3665), .Y(N152) );
  MXI4X1 U4203 ( .A(\block[0][0][22] ), .B(\block[1][0][22] ), .C(
        \block[2][0][22] ), .D(\block[3][0][22] ), .S0(n3619), .S1(n3651), .Y(
        n3550) );
  MXI4X1 U4204 ( .A(\block[4][0][22] ), .B(\block[5][0][22] ), .C(
        \block[6][0][22] ), .D(\block[7][0][22] ), .S0(n3619), .S1(n3651), .Y(
        n3551) );
  MXI2X1 U4205 ( .A(n3548), .B(n3549), .S0(n3665), .Y(N151) );
  MXI4X1 U4206 ( .A(\block[0][0][23] ), .B(\block[1][0][23] ), .C(
        \block[2][0][23] ), .D(\block[3][0][23] ), .S0(n3619), .S1(n3651), .Y(
        n3548) );
  MXI4X1 U4207 ( .A(\block[4][0][23] ), .B(\block[5][0][23] ), .C(
        \block[6][0][23] ), .D(\block[7][0][23] ), .S0(n3619), .S1(n3651), .Y(
        n3549) );
  MXI2X1 U4208 ( .A(n3546), .B(n3547), .S0(n3664), .Y(N150) );
  MXI4X1 U4209 ( .A(\block[0][0][24] ), .B(\block[1][0][24] ), .C(
        \block[2][0][24] ), .D(\block[3][0][24] ), .S0(n3619), .S1(n3650), .Y(
        n3546) );
  MXI4X1 U4210 ( .A(\block[4][0][24] ), .B(\block[5][0][24] ), .C(
        \block[6][0][24] ), .D(\block[7][0][24] ), .S0(n3619), .S1(n3650), .Y(
        n3547) );
  MXI2X1 U4211 ( .A(n3544), .B(n3545), .S0(n3664), .Y(N149) );
  MXI4X1 U4212 ( .A(\block[0][0][25] ), .B(\block[1][0][25] ), .C(
        \block[2][0][25] ), .D(\block[3][0][25] ), .S0(n3619), .S1(n3650), .Y(
        n3544) );
  MXI4X1 U4213 ( .A(\block[4][0][25] ), .B(\block[5][0][25] ), .C(
        \block[6][0][25] ), .D(\block[7][0][25] ), .S0(n3619), .S1(n3650), .Y(
        n3545) );
  MXI2X1 U4214 ( .A(n3542), .B(n3543), .S0(n3664), .Y(N148) );
  MXI4X1 U4215 ( .A(\block[0][0][26] ), .B(\block[1][0][26] ), .C(
        \block[2][0][26] ), .D(\block[3][0][26] ), .S0(n3620), .S1(n3650), .Y(
        n3542) );
  MXI4X1 U4216 ( .A(\block[4][0][26] ), .B(\block[5][0][26] ), .C(
        \block[6][0][26] ), .D(\block[7][0][26] ), .S0(n3608), .S1(n3650), .Y(
        n3543) );
  MXI2X1 U4217 ( .A(n3540), .B(n3541), .S0(n3664), .Y(N147) );
  MXI4X1 U4218 ( .A(\block[0][0][27] ), .B(\block[1][0][27] ), .C(
        \block[2][0][27] ), .D(\block[3][0][27] ), .S0(n3621), .S1(n3650), .Y(
        n3540) );
  MXI4X1 U4219 ( .A(\block[4][0][27] ), .B(\block[5][0][27] ), .C(
        \block[6][0][27] ), .D(\block[7][0][27] ), .S0(n3609), .S1(n3650), .Y(
        n3541) );
  MXI2X1 U4220 ( .A(n3538), .B(n3539), .S0(n3664), .Y(N146) );
  MXI4X1 U4221 ( .A(\block[0][0][28] ), .B(\block[1][0][28] ), .C(
        \block[2][0][28] ), .D(\block[3][0][28] ), .S0(n3620), .S1(n3650), .Y(
        n3538) );
  MXI4X1 U4222 ( .A(\block[4][0][28] ), .B(\block[5][0][28] ), .C(
        \block[6][0][28] ), .D(\block[7][0][28] ), .S0(n3614), .S1(n3650), .Y(
        n3539) );
  MXI2X1 U4223 ( .A(n3536), .B(n3537), .S0(n3664), .Y(N145) );
  MXI4X1 U4224 ( .A(\block[0][0][29] ), .B(\block[1][0][29] ), .C(
        \block[2][0][29] ), .D(\block[3][0][29] ), .S0(n3621), .S1(n3650), .Y(
        n3536) );
  MXI4X1 U4225 ( .A(\block[4][0][29] ), .B(\block[5][0][29] ), .C(
        \block[6][0][29] ), .D(\block[7][0][29] ), .S0(n3613), .S1(n3650), .Y(
        n3537) );
  MXI2X1 U4226 ( .A(n3534), .B(n3535), .S0(n3664), .Y(N144) );
  MXI4X1 U4227 ( .A(\block[0][0][30] ), .B(\block[1][0][30] ), .C(
        \block[2][0][30] ), .D(\block[3][0][30] ), .S0(n3612), .S1(n3649), .Y(
        n3534) );
  MXI4X1 U4228 ( .A(\block[4][0][30] ), .B(\block[5][0][30] ), .C(
        \block[6][0][30] ), .D(\block[7][0][30] ), .S0(n3619), .S1(n3649), .Y(
        n3535) );
  MXI2X1 U4229 ( .A(n3532), .B(n3533), .S0(n3664), .Y(N143) );
  MXI4X1 U4230 ( .A(\block[0][0][31] ), .B(\block[1][0][31] ), .C(
        \block[2][0][31] ), .D(\block[3][0][31] ), .S0(n3617), .S1(n3649), .Y(
        n3532) );
  MXI4X1 U4231 ( .A(\block[4][0][31] ), .B(\block[5][0][31] ), .C(
        \block[6][0][31] ), .D(\block[7][0][31] ), .S0(n3610), .S1(n3649), .Y(
        n3533) );
  MXI2X1 U4232 ( .A(n3402), .B(n3403), .S0(n3660), .Y(N78) );
  MXI4X1 U4233 ( .A(\block[0][3][0] ), .B(\block[1][3][0] ), .C(
        \block[2][3][0] ), .D(\block[3][3][0] ), .S0(n3611), .S1(n3639), .Y(
        n3402) );
  MXI4X1 U4234 ( .A(\block[4][3][0] ), .B(\block[5][3][0] ), .C(
        \block[6][3][0] ), .D(\block[7][3][0] ), .S0(n3611), .S1(n3639), .Y(
        n3403) );
  MXI2X1 U4235 ( .A(n3400), .B(n3401), .S0(n3660), .Y(N77) );
  MXI4X1 U4236 ( .A(\block[0][3][1] ), .B(\block[1][3][1] ), .C(
        \block[2][3][1] ), .D(\block[3][3][1] ), .S0(n3611), .S1(n3639), .Y(
        n3400) );
  MXI4X1 U4237 ( .A(\block[4][3][1] ), .B(\block[5][3][1] ), .C(
        \block[6][3][1] ), .D(\block[7][3][1] ), .S0(n3610), .S1(n3639), .Y(
        n3401) );
  MXI2X1 U4238 ( .A(n3398), .B(n3399), .S0(n3660), .Y(N76) );
  MXI4X1 U4239 ( .A(\block[0][3][2] ), .B(\block[1][3][2] ), .C(
        \block[2][3][2] ), .D(\block[3][3][2] ), .S0(n3610), .S1(n3639), .Y(
        n3398) );
  MXI4X1 U4240 ( .A(\block[4][3][2] ), .B(\block[5][3][2] ), .C(
        \block[6][3][2] ), .D(\block[7][3][2] ), .S0(n3610), .S1(n3639), .Y(
        n3399) );
  MXI2X1 U4241 ( .A(n3396), .B(n3397), .S0(n3660), .Y(N75) );
  MXI4X1 U4242 ( .A(\block[0][3][3] ), .B(\block[1][3][3] ), .C(
        \block[2][3][3] ), .D(\block[3][3][3] ), .S0(n3610), .S1(n3639), .Y(
        n3396) );
  MXI4X1 U4243 ( .A(\block[4][3][3] ), .B(\block[5][3][3] ), .C(
        \block[6][3][3] ), .D(\block[7][3][3] ), .S0(n3610), .S1(n3639), .Y(
        n3397) );
  MXI2X1 U4244 ( .A(n3394), .B(n3395), .S0(n3660), .Y(N74) );
  MXI4X1 U4245 ( .A(\block[0][3][4] ), .B(\block[1][3][4] ), .C(
        \block[2][3][4] ), .D(\block[3][3][4] ), .S0(n3610), .S1(n3639), .Y(
        n3394) );
  MXI4X1 U4246 ( .A(\block[4][3][4] ), .B(\block[5][3][4] ), .C(
        \block[6][3][4] ), .D(\block[7][3][4] ), .S0(n3610), .S1(n3639), .Y(
        n3395) );
  MXI2X1 U4247 ( .A(n3392), .B(n3393), .S0(n3660), .Y(N73) );
  MXI4X1 U4248 ( .A(\block[0][3][5] ), .B(\block[1][3][5] ), .C(
        \block[2][3][5] ), .D(\block[3][3][5] ), .S0(n3610), .S1(n3639), .Y(
        n3392) );
  MXI4X1 U4249 ( .A(\block[4][3][5] ), .B(\block[5][3][5] ), .C(
        \block[6][3][5] ), .D(\block[7][3][5] ), .S0(n3610), .S1(n3639), .Y(
        n3393) );
  MXI2X1 U4250 ( .A(n3390), .B(n3391), .S0(n3660), .Y(N72) );
  MXI4X1 U4251 ( .A(\block[0][3][6] ), .B(\block[1][3][6] ), .C(
        \block[2][3][6] ), .D(\block[3][3][6] ), .S0(n3610), .S1(n3638), .Y(
        n3390) );
  MXI4X1 U4252 ( .A(\block[4][3][6] ), .B(\block[5][3][6] ), .C(
        \block[6][3][6] ), .D(\block[7][3][6] ), .S0(n3610), .S1(n3638), .Y(
        n3391) );
  MXI2X1 U4253 ( .A(n3388), .B(n3389), .S0(n3660), .Y(N71) );
  MXI4X1 U4254 ( .A(\block[0][3][7] ), .B(\block[1][3][7] ), .C(
        \block[2][3][7] ), .D(\block[3][3][7] ), .S0(n3610), .S1(n3638), .Y(
        n3388) );
  MXI4X1 U4255 ( .A(\block[4][3][7] ), .B(\block[5][3][7] ), .C(
        \block[6][3][7] ), .D(\block[7][3][7] ), .S0(n3610), .S1(n3638), .Y(
        n3389) );
  MXI2X1 U4256 ( .A(n3386), .B(n3387), .S0(n3660), .Y(N70) );
  MXI4X1 U4257 ( .A(\block[0][3][8] ), .B(\block[1][3][8] ), .C(
        \block[2][3][8] ), .D(\block[3][3][8] ), .S0(n3609), .S1(n3638), .Y(
        n3386) );
  MXI4X1 U4258 ( .A(\block[4][3][8] ), .B(\block[5][3][8] ), .C(
        \block[6][3][8] ), .D(\block[7][3][8] ), .S0(n3609), .S1(n3638), .Y(
        n3387) );
  MXI2X1 U4259 ( .A(n3384), .B(n3385), .S0(n3660), .Y(N69) );
  MXI4X1 U4260 ( .A(\block[0][3][9] ), .B(\block[1][3][9] ), .C(
        \block[2][3][9] ), .D(\block[3][3][9] ), .S0(n3609), .S1(n3638), .Y(
        n3384) );
  MXI4X1 U4261 ( .A(\block[4][3][9] ), .B(\block[5][3][9] ), .C(
        \block[6][3][9] ), .D(\block[7][3][9] ), .S0(n3609), .S1(n3638), .Y(
        n3385) );
  MXI2X1 U4262 ( .A(n3382), .B(n3383), .S0(n3660), .Y(N68) );
  MXI4X1 U4263 ( .A(\block[0][3][10] ), .B(\block[1][3][10] ), .C(
        \block[2][3][10] ), .D(\block[3][3][10] ), .S0(n3609), .S1(n3638), .Y(
        n3382) );
  MXI4X1 U4264 ( .A(\block[4][3][10] ), .B(\block[5][3][10] ), .C(
        \block[6][3][10] ), .D(\block[7][3][10] ), .S0(n3609), .S1(n3638), .Y(
        n3383) );
  MXI2X1 U4265 ( .A(n3380), .B(n3381), .S0(n3660), .Y(N67) );
  MXI4X1 U4266 ( .A(\block[0][3][11] ), .B(\block[1][3][11] ), .C(
        \block[2][3][11] ), .D(\block[3][3][11] ), .S0(n3609), .S1(n3638), .Y(
        n3380) );
  MXI4X1 U4267 ( .A(\block[4][3][11] ), .B(\block[5][3][11] ), .C(
        \block[6][3][11] ), .D(\block[7][3][11] ), .S0(n3609), .S1(n3638), .Y(
        n3381) );
  MXI2X1 U4268 ( .A(n3378), .B(n3379), .S0(n3661), .Y(N66) );
  MXI4X1 U4269 ( .A(\block[0][3][12] ), .B(\block[1][3][12] ), .C(
        \block[2][3][12] ), .D(\block[3][3][12] ), .S0(n3609), .S1(n3637), .Y(
        n3378) );
  MXI4X1 U4270 ( .A(\block[4][3][12] ), .B(\block[5][3][12] ), .C(
        \block[6][3][12] ), .D(\block[7][3][12] ), .S0(n3609), .S1(n3637), .Y(
        n3379) );
  MXI2X1 U4271 ( .A(n3376), .B(n3377), .S0(n3658), .Y(N65) );
  MXI4X1 U4272 ( .A(\block[0][3][13] ), .B(\block[1][3][13] ), .C(
        \block[2][3][13] ), .D(\block[3][3][13] ), .S0(n3609), .S1(n3637), .Y(
        n3376) );
  MXI4X1 U4273 ( .A(\block[4][3][13] ), .B(\block[5][3][13] ), .C(
        \block[6][3][13] ), .D(\block[7][3][13] ), .S0(n3609), .S1(n3637), .Y(
        n3377) );
  MXI2X1 U4274 ( .A(n3374), .B(n3375), .S0(n3658), .Y(N64) );
  MXI4X1 U4275 ( .A(\block[0][3][14] ), .B(\block[1][3][14] ), .C(
        \block[2][3][14] ), .D(\block[3][3][14] ), .S0(n3609), .S1(n3637), .Y(
        n3374) );
  MXI4X1 U4276 ( .A(\block[4][3][14] ), .B(\block[5][3][14] ), .C(
        \block[6][3][14] ), .D(\block[7][3][14] ), .S0(n3608), .S1(n3637), .Y(
        n3375) );
  MXI2X1 U4277 ( .A(n3372), .B(n3373), .S0(n3658), .Y(N63) );
  MXI4X1 U4278 ( .A(\block[0][3][15] ), .B(\block[1][3][15] ), .C(
        \block[2][3][15] ), .D(\block[3][3][15] ), .S0(n3608), .S1(n3637), .Y(
        n3372) );
  MXI4X1 U4279 ( .A(\block[4][3][15] ), .B(\block[5][3][15] ), .C(
        \block[6][3][15] ), .D(\block[7][3][15] ), .S0(n3608), .S1(n3637), .Y(
        n3373) );
  MXI2X1 U4280 ( .A(n3370), .B(n3371), .S0(n3658), .Y(N62) );
  MXI4X1 U4281 ( .A(\block[0][3][16] ), .B(\block[1][3][16] ), .C(
        \block[2][3][16] ), .D(\block[3][3][16] ), .S0(n3608), .S1(n3637), .Y(
        n3370) );
  MXI4X1 U4282 ( .A(\block[4][3][16] ), .B(\block[5][3][16] ), .C(
        \block[6][3][16] ), .D(\block[7][3][16] ), .S0(n3608), .S1(n3637), .Y(
        n3371) );
  MXI2X1 U4283 ( .A(n3368), .B(n3369), .S0(n3662), .Y(N61) );
  MXI4X1 U4284 ( .A(\block[0][3][17] ), .B(\block[1][3][17] ), .C(
        \block[2][3][17] ), .D(\block[3][3][17] ), .S0(n3608), .S1(n3637), .Y(
        n3368) );
  MXI4X1 U4285 ( .A(\block[4][3][17] ), .B(\block[5][3][17] ), .C(
        \block[6][3][17] ), .D(\block[7][3][17] ), .S0(n3608), .S1(n3637), .Y(
        n3369) );
  MXI2X1 U4286 ( .A(n3366), .B(n3367), .S0(n3658), .Y(N60) );
  MXI4X1 U4287 ( .A(\block[0][3][18] ), .B(\block[1][3][18] ), .C(
        \block[2][3][18] ), .D(\block[3][3][18] ), .S0(n3608), .S1(n3636), .Y(
        n3366) );
  MXI4X1 U4288 ( .A(\block[4][3][18] ), .B(\block[5][3][18] ), .C(
        \block[6][3][18] ), .D(\block[7][3][18] ), .S0(n3608), .S1(n3636), .Y(
        n3367) );
  MXI2X1 U4289 ( .A(n3364), .B(n3365), .S0(n3662), .Y(N59) );
  MXI4X1 U4290 ( .A(\block[0][3][19] ), .B(\block[1][3][19] ), .C(
        \block[2][3][19] ), .D(\block[3][3][19] ), .S0(n3608), .S1(n3636), .Y(
        n3364) );
  MXI4X1 U4291 ( .A(\block[4][3][19] ), .B(\block[5][3][19] ), .C(
        \block[6][3][19] ), .D(\block[7][3][19] ), .S0(n3608), .S1(n3636), .Y(
        n3365) );
  MXI2X1 U4292 ( .A(n3362), .B(n3363), .S0(n3658), .Y(N58) );
  MXI4X1 U4293 ( .A(\block[0][3][20] ), .B(\block[1][3][20] ), .C(
        \block[2][3][20] ), .D(\block[3][3][20] ), .S0(n3608), .S1(n3636), .Y(
        n3362) );
  MXI4X1 U4294 ( .A(\block[4][3][20] ), .B(\block[5][3][20] ), .C(
        \block[6][3][20] ), .D(\block[7][3][20] ), .S0(n3608), .S1(n3636), .Y(
        n3363) );
  MXI2X1 U4295 ( .A(n3360), .B(n3361), .S0(n3658), .Y(N57) );
  MXI4X1 U4296 ( .A(\block[0][3][21] ), .B(\block[1][3][21] ), .C(
        \block[2][3][21] ), .D(\block[3][3][21] ), .S0(n3607), .S1(n3636), .Y(
        n3360) );
  MXI4X1 U4297 ( .A(\block[4][3][21] ), .B(\block[5][3][21] ), .C(
        \block[6][3][21] ), .D(\block[7][3][21] ), .S0(n3607), .S1(n3636), .Y(
        n3361) );
  MXI2X1 U4298 ( .A(n3358), .B(n3359), .S0(n3660), .Y(N56) );
  MXI4X1 U4299 ( .A(\block[0][3][22] ), .B(\block[1][3][22] ), .C(
        \block[2][3][22] ), .D(\block[3][3][22] ), .S0(n3607), .S1(n3636), .Y(
        n3358) );
  MXI4X1 U4300 ( .A(\block[4][3][22] ), .B(\block[5][3][22] ), .C(
        \block[6][3][22] ), .D(\block[7][3][22] ), .S0(n3607), .S1(n3636), .Y(
        n3359) );
  MXI2X1 U4301 ( .A(n3356), .B(n3357), .S0(n3658), .Y(N55) );
  MXI4X1 U4302 ( .A(\block[0][3][23] ), .B(\block[1][3][23] ), .C(
        \block[2][3][23] ), .D(\block[3][3][23] ), .S0(n3607), .S1(n3636), .Y(
        n3356) );
  MXI4X1 U4303 ( .A(\block[4][3][23] ), .B(\block[5][3][23] ), .C(
        \block[6][3][23] ), .D(\block[7][3][23] ), .S0(n3607), .S1(n3636), .Y(
        n3357) );
  MXI4X1 U4304 ( .A(\block[0][3][24] ), .B(\block[1][3][24] ), .C(
        \block[2][3][24] ), .D(\block[3][3][24] ), .S0(n3607), .S1(n3635), .Y(
        n3354) );
  MXI4X1 U4305 ( .A(\block[4][3][24] ), .B(\block[5][3][24] ), .C(
        \block[6][3][24] ), .D(\block[7][3][24] ), .S0(n3607), .S1(n3635), .Y(
        n3355) );
  MXI4X1 U4306 ( .A(\block[0][3][25] ), .B(\block[1][3][25] ), .C(
        \block[2][3][25] ), .D(\block[3][3][25] ), .S0(n3607), .S1(n3635), .Y(
        n3352) );
  MXI4X1 U4307 ( .A(\block[4][3][25] ), .B(\block[5][3][25] ), .C(
        \block[6][3][25] ), .D(\block[7][3][25] ), .S0(n3607), .S1(n3635), .Y(
        n3353) );
  MXI4X1 U4308 ( .A(\block[0][3][26] ), .B(\block[1][3][26] ), .C(
        \block[2][3][26] ), .D(\block[3][3][26] ), .S0(n3607), .S1(n3635), .Y(
        n3350) );
  MXI4X1 U4309 ( .A(\block[4][3][26] ), .B(\block[5][3][26] ), .C(
        \block[6][3][26] ), .D(\block[7][3][26] ), .S0(n3607), .S1(n3635), .Y(
        n3351) );
  MXI4X1 U4310 ( .A(\block[0][3][27] ), .B(\block[1][3][27] ), .C(
        \block[2][3][27] ), .D(\block[3][3][27] ), .S0(n3607), .S1(n3635), .Y(
        n3348) );
  MXI2X1 U4311 ( .A(n3530), .B(n3531), .S0(n3664), .Y(N142) );
  MXI4X1 U4312 ( .A(\block[0][1][0] ), .B(\block[1][1][0] ), .C(
        \block[2][1][0] ), .D(\block[3][1][0] ), .S0(n3617), .S1(n3649), .Y(
        n3530) );
  MXI4X1 U4313 ( .A(\block[4][1][0] ), .B(\block[5][1][0] ), .C(
        \block[6][1][0] ), .D(\block[7][1][0] ), .S0(n3618), .S1(n3649), .Y(
        n3531) );
  MXI2X1 U4314 ( .A(n3528), .B(n3529), .S0(n3664), .Y(N141) );
  MXI4X1 U4315 ( .A(\block[0][1][1] ), .B(\block[1][1][1] ), .C(
        \block[2][1][1] ), .D(\block[3][1][1] ), .S0(n3618), .S1(n3649), .Y(
        n3528) );
  MXI4X1 U4316 ( .A(\block[4][1][1] ), .B(\block[5][1][1] ), .C(
        \block[6][1][1] ), .D(\block[7][1][1] ), .S0(n3618), .S1(n3649), .Y(
        n3529) );
  MXI2X1 U4317 ( .A(n3526), .B(n3527), .S0(n3664), .Y(N140) );
  MXI4X1 U4318 ( .A(\block[0][1][2] ), .B(\block[1][1][2] ), .C(
        \block[2][1][2] ), .D(\block[3][1][2] ), .S0(n3618), .S1(n3649), .Y(
        n3526) );
  MXI4X1 U4319 ( .A(\block[4][1][2] ), .B(\block[5][1][2] ), .C(
        \block[6][1][2] ), .D(\block[7][1][2] ), .S0(n3618), .S1(n3649), .Y(
        n3527) );
  MXI2X1 U4320 ( .A(n3524), .B(n3525), .S0(n3664), .Y(N139) );
  MXI4X1 U4321 ( .A(\block[0][1][3] ), .B(\block[1][1][3] ), .C(
        \block[2][1][3] ), .D(\block[3][1][3] ), .S0(n3618), .S1(n3649), .Y(
        n3524) );
  MXI4X1 U4322 ( .A(\block[4][1][3] ), .B(\block[5][1][3] ), .C(
        \block[6][1][3] ), .D(\block[7][1][3] ), .S0(n3618), .S1(n3649), .Y(
        n3525) );
  MXI2X1 U4323 ( .A(n3522), .B(n3523), .S0(n3663), .Y(N138) );
  MXI4X1 U4324 ( .A(\block[0][1][4] ), .B(\block[1][1][4] ), .C(
        \block[2][1][4] ), .D(\block[3][1][4] ), .S0(n3618), .S1(n3648), .Y(
        n3522) );
  MXI4X1 U4325 ( .A(\block[4][1][4] ), .B(\block[5][1][4] ), .C(
        \block[6][1][4] ), .D(\block[7][1][4] ), .S0(n3618), .S1(n3648), .Y(
        n3523) );
  MXI2X1 U4326 ( .A(n3520), .B(n3521), .S0(n3663), .Y(N137) );
  MXI4X1 U4327 ( .A(\block[0][1][5] ), .B(\block[1][1][5] ), .C(
        \block[2][1][5] ), .D(\block[3][1][5] ), .S0(n3618), .S1(n3648), .Y(
        n3520) );
  MXI4X1 U4328 ( .A(\block[4][1][5] ), .B(\block[5][1][5] ), .C(
        \block[6][1][5] ), .D(\block[7][1][5] ), .S0(n3618), .S1(n3648), .Y(
        n3521) );
  MXI2X1 U4329 ( .A(n3518), .B(n3519), .S0(n3663), .Y(N136) );
  MXI4X1 U4330 ( .A(\block[0][1][6] ), .B(\block[1][1][6] ), .C(
        \block[2][1][6] ), .D(\block[3][1][6] ), .S0(n3618), .S1(n3648), .Y(
        n3518) );
  MXI4X1 U4331 ( .A(\block[4][1][6] ), .B(\block[5][1][6] ), .C(
        \block[6][1][6] ), .D(\block[7][1][6] ), .S0(n3618), .S1(n3648), .Y(
        n3519) );
  MXI2X1 U4332 ( .A(n3516), .B(n3517), .S0(n3663), .Y(N135) );
  MXI4X1 U4333 ( .A(\block[0][1][7] ), .B(\block[1][1][7] ), .C(
        \block[2][1][7] ), .D(\block[3][1][7] ), .S0(n3617), .S1(n3648), .Y(
        n3516) );
  MXI4X1 U4334 ( .A(\block[4][1][7] ), .B(\block[5][1][7] ), .C(
        \block[6][1][7] ), .D(\block[7][1][7] ), .S0(n3617), .S1(n3648), .Y(
        n3517) );
  MXI2X1 U4335 ( .A(n3514), .B(n3515), .S0(n3663), .Y(N134) );
  MXI4X1 U4336 ( .A(\block[0][1][8] ), .B(\block[1][1][8] ), .C(
        \block[2][1][8] ), .D(\block[3][1][8] ), .S0(n3617), .S1(n3648), .Y(
        n3514) );
  MXI4X1 U4337 ( .A(\block[4][1][8] ), .B(\block[5][1][8] ), .C(
        \block[6][1][8] ), .D(\block[7][1][8] ), .S0(n3617), .S1(n3648), .Y(
        n3515) );
  MXI2X1 U4338 ( .A(n3512), .B(n3513), .S0(n3663), .Y(N133) );
  MXI4X1 U4339 ( .A(\block[0][1][9] ), .B(\block[1][1][9] ), .C(
        \block[2][1][9] ), .D(\block[3][1][9] ), .S0(n3617), .S1(n3648), .Y(
        n3512) );
  MXI4X1 U4340 ( .A(\block[4][1][9] ), .B(\block[5][1][9] ), .C(
        \block[6][1][9] ), .D(\block[7][1][9] ), .S0(n3617), .S1(n3648), .Y(
        n3513) );
  MXI2X1 U4341 ( .A(n3510), .B(n3511), .S0(n3663), .Y(N132) );
  MXI4X1 U4342 ( .A(\block[0][1][10] ), .B(\block[1][1][10] ), .C(
        \block[2][1][10] ), .D(\block[3][1][10] ), .S0(n3617), .S1(n3647), .Y(
        n3510) );
  MXI4X1 U4343 ( .A(\block[4][1][10] ), .B(\block[5][1][10] ), .C(
        \block[6][1][10] ), .D(\block[7][1][10] ), .S0(n3617), .S1(n3647), .Y(
        n3511) );
  MXI2X1 U4344 ( .A(n3508), .B(n3509), .S0(n3663), .Y(N131) );
  MXI4X1 U4345 ( .A(\block[0][1][11] ), .B(\block[1][1][11] ), .C(
        \block[2][1][11] ), .D(\block[3][1][11] ), .S0(n3617), .S1(n3647), .Y(
        n3508) );
  MXI4X1 U4346 ( .A(\block[4][1][11] ), .B(\block[5][1][11] ), .C(
        \block[6][1][11] ), .D(\block[7][1][11] ), .S0(n3617), .S1(n3647), .Y(
        n3509) );
  MXI2X1 U4347 ( .A(n3506), .B(n3507), .S0(n3663), .Y(N130) );
  MXI4X1 U4348 ( .A(\block[0][1][12] ), .B(\block[1][1][12] ), .C(
        \block[2][1][12] ), .D(\block[3][1][12] ), .S0(n3617), .S1(n3647), .Y(
        n3506) );
  MXI4X1 U4349 ( .A(\block[4][1][12] ), .B(\block[5][1][12] ), .C(
        \block[6][1][12] ), .D(\block[7][1][12] ), .S0(n3617), .S1(n3647), .Y(
        n3507) );
  MXI2X1 U4350 ( .A(n3504), .B(n3505), .S0(n3663), .Y(N129) );
  MXI4X1 U4351 ( .A(\block[0][1][13] ), .B(\block[1][1][13] ), .C(
        \block[2][1][13] ), .D(\block[3][1][13] ), .S0(n3617), .S1(n3647), .Y(
        n3504) );
  MXI4X1 U4352 ( .A(\block[4][1][13] ), .B(\block[5][1][13] ), .C(
        \block[6][1][13] ), .D(\block[7][1][13] ), .S0(n3618), .S1(n3647), .Y(
        n3505) );
  MXI2X1 U4353 ( .A(n3502), .B(n3503), .S0(n3663), .Y(N128) );
  MXI4X1 U4354 ( .A(\block[0][1][14] ), .B(\block[1][1][14] ), .C(
        \block[2][1][14] ), .D(\block[3][1][14] ), .S0(n3610), .S1(n3647), .Y(
        n3502) );
  MXI4X1 U4355 ( .A(\block[4][1][14] ), .B(\block[5][1][14] ), .C(
        \block[6][1][14] ), .D(\block[7][1][14] ), .S0(n3610), .S1(n3647), .Y(
        n3503) );
  MXI2X1 U4356 ( .A(n3500), .B(n3501), .S0(n3663), .Y(N127) );
  MXI4X1 U4357 ( .A(\block[0][1][15] ), .B(\block[1][1][15] ), .C(
        \block[2][1][15] ), .D(\block[3][1][15] ), .S0(n3620), .S1(n3647), .Y(
        n3500) );
  MXI4X1 U4358 ( .A(\block[4][1][15] ), .B(\block[5][1][15] ), .C(
        \block[6][1][15] ), .D(\block[7][1][15] ), .S0(n3611), .S1(n3647), .Y(
        n3501) );
  MXI2X1 U4359 ( .A(n3498), .B(n3499), .S0(n3663), .Y(N126) );
  MXI4X1 U4360 ( .A(\block[0][1][16] ), .B(\block[1][1][16] ), .C(
        \block[2][1][16] ), .D(\block[3][1][16] ), .S0(n3613), .S1(n3646), .Y(
        n3498) );
  MXI4X1 U4361 ( .A(\block[4][1][16] ), .B(\block[5][1][16] ), .C(
        \block[6][1][16] ), .D(\block[7][1][16] ), .S0(n3613), .S1(n3646), .Y(
        n3499) );
  MXI2X1 U4362 ( .A(n3496), .B(n3497), .S0(n3663), .Y(N125) );
  MXI4X1 U4363 ( .A(\block[0][1][17] ), .B(\block[1][1][17] ), .C(
        \block[2][1][17] ), .D(\block[3][1][17] ), .S0(n3619), .S1(n3646), .Y(
        n3496) );
  MXI4X1 U4364 ( .A(\block[4][1][17] ), .B(\block[5][1][17] ), .C(
        \block[6][1][17] ), .D(\block[7][1][17] ), .S0(n3619), .S1(n3646), .Y(
        n3497) );
  MXI2X1 U4365 ( .A(n3494), .B(n3495), .S0(n3663), .Y(N124) );
  MXI4X1 U4366 ( .A(\block[0][1][18] ), .B(\block[1][1][18] ), .C(
        \block[2][1][18] ), .D(\block[3][1][18] ), .S0(n3612), .S1(n3646), .Y(
        n3494) );
  MXI4X1 U4367 ( .A(\block[4][1][18] ), .B(\block[5][1][18] ), .C(
        \block[6][1][18] ), .D(\block[7][1][18] ), .S0(n3612), .S1(n3646), .Y(
        n3495) );
  MXI2X1 U4368 ( .A(n3492), .B(n3493), .S0(n3664), .Y(N123) );
  MXI4X1 U4369 ( .A(\block[0][1][19] ), .B(\block[1][1][19] ), .C(
        \block[2][1][19] ), .D(\block[3][1][19] ), .S0(n3618), .S1(n3646), .Y(
        n3492) );
  MXI4X1 U4370 ( .A(\block[4][1][19] ), .B(\block[5][1][19] ), .C(
        \block[6][1][19] ), .D(\block[7][1][19] ), .S0(n3618), .S1(n3646), .Y(
        n3493) );
  MXI2X1 U4371 ( .A(n3490), .B(n3491), .S0(n3666), .Y(N122) );
  MXI4X1 U4372 ( .A(\block[0][1][20] ), .B(\block[1][1][20] ), .C(
        \block[2][1][20] ), .D(\block[3][1][20] ), .S0(n3616), .S1(n3646), .Y(
        n3490) );
  MXI4X1 U4373 ( .A(\block[4][1][20] ), .B(\block[5][1][20] ), .C(
        \block[6][1][20] ), .D(\block[7][1][20] ), .S0(n3616), .S1(n3646), .Y(
        n3491) );
  MXI2X1 U4374 ( .A(n3488), .B(n3489), .S0(n3665), .Y(N121) );
  MXI4X1 U4375 ( .A(\block[0][1][21] ), .B(\block[1][1][21] ), .C(
        \block[2][1][21] ), .D(\block[3][1][21] ), .S0(n3616), .S1(n3646), .Y(
        n3488) );
  MXI4X1 U4376 ( .A(\block[4][1][21] ), .B(\block[5][1][21] ), .C(
        \block[6][1][21] ), .D(\block[7][1][21] ), .S0(n3616), .S1(n3646), .Y(
        n3489) );
  MXI2X1 U4377 ( .A(n3486), .B(n3487), .S0(n3664), .Y(N120) );
  MXI4X1 U4378 ( .A(\block[0][1][22] ), .B(\block[1][1][22] ), .C(
        \block[2][1][22] ), .D(\block[3][1][22] ), .S0(n3616), .S1(n3653), .Y(
        n3486) );
  MXI4X1 U4379 ( .A(\block[4][1][22] ), .B(\block[5][1][22] ), .C(
        \block[6][1][22] ), .D(\block[7][1][22] ), .S0(n3616), .S1(n3653), .Y(
        n3487) );
  MXI2X1 U4380 ( .A(n3484), .B(n3485), .S0(n3663), .Y(N119) );
  MXI4X1 U4381 ( .A(\block[0][1][23] ), .B(\block[1][1][23] ), .C(
        \block[2][1][23] ), .D(\block[3][1][23] ), .S0(n3616), .S1(n3654), .Y(
        n3484) );
  MXI4X1 U4382 ( .A(\block[4][1][23] ), .B(\block[5][1][23] ), .C(
        \block[6][1][23] ), .D(\block[7][1][23] ), .S0(n3616), .S1(n3654), .Y(
        n3485) );
  MXI2X1 U4383 ( .A(n3482), .B(n3483), .S0(n3664), .Y(N118) );
  MXI4X1 U4384 ( .A(\block[0][1][24] ), .B(\block[1][1][24] ), .C(
        \block[2][1][24] ), .D(\block[3][1][24] ), .S0(n3616), .S1(n3646), .Y(
        n3482) );
  MXI4X1 U4385 ( .A(\block[4][1][24] ), .B(\block[5][1][24] ), .C(
        \block[6][1][24] ), .D(\block[7][1][24] ), .S0(n3616), .S1(n3646), .Y(
        n3483) );
  MXI2X1 U4386 ( .A(n3480), .B(n3481), .S0(n3664), .Y(N117) );
  MXI4X1 U4387 ( .A(\block[0][1][25] ), .B(\block[1][1][25] ), .C(
        \block[2][1][25] ), .D(\block[3][1][25] ), .S0(n3616), .S1(n3652), .Y(
        n3480) );
  MXI4X1 U4388 ( .A(\block[4][1][25] ), .B(\block[5][1][25] ), .C(
        \block[6][1][25] ), .D(\block[7][1][25] ), .S0(n3616), .S1(n3652), .Y(
        n3481) );
  MXI2X1 U4389 ( .A(n3478), .B(n3479), .S0(n3663), .Y(N116) );
  MXI4X1 U4390 ( .A(\block[0][1][26] ), .B(\block[1][1][26] ), .C(
        \block[2][1][26] ), .D(\block[3][1][26] ), .S0(n3616), .S1(n3651), .Y(
        n3478) );
  MXI4X1 U4391 ( .A(\block[4][1][26] ), .B(\block[5][1][26] ), .C(
        \block[6][1][26] ), .D(\block[7][1][26] ), .S0(n3616), .S1(n3651), .Y(
        n3479) );
  MXI2X1 U4392 ( .A(n3476), .B(n3477), .S0(n3664), .Y(N115) );
  MXI4X1 U4393 ( .A(\block[0][1][27] ), .B(\block[1][1][27] ), .C(
        \block[2][1][27] ), .D(\block[3][1][27] ), .S0(n3609), .S1(n3641), .Y(
        n3476) );
  MXI4X1 U4394 ( .A(\block[4][1][27] ), .B(\block[5][1][27] ), .C(
        \block[6][1][27] ), .D(\block[7][1][27] ), .S0(n3608), .S1(n3641), .Y(
        n3477) );
  MXI2X1 U4395 ( .A(n3474), .B(n3475), .S0(n3661), .Y(N114) );
  MXI4X1 U4396 ( .A(\block[0][1][28] ), .B(\block[1][1][28] ), .C(
        \block[2][1][28] ), .D(\block[3][1][28] ), .S0(n3614), .S1(n3645), .Y(
        n3474) );
  MXI4X1 U4397 ( .A(\block[4][1][28] ), .B(\block[5][1][28] ), .C(
        \block[6][1][28] ), .D(\block[7][1][28] ), .S0(n3614), .S1(n3645), .Y(
        n3475) );
  MXI2X1 U4398 ( .A(n3472), .B(n3473), .S0(n3660), .Y(N113) );
  MXI4X1 U4399 ( .A(\block[0][1][29] ), .B(\block[1][1][29] ), .C(
        \block[2][1][29] ), .D(\block[3][1][29] ), .S0(n3615), .S1(n3645), .Y(
        n3472) );
  MXI4X1 U4400 ( .A(\block[4][1][29] ), .B(\block[5][1][29] ), .C(
        \block[6][1][29] ), .D(\block[7][1][29] ), .S0(n3615), .S1(n3645), .Y(
        n3473) );
  MXI2X1 U4401 ( .A(n3470), .B(n3471), .S0(n3660), .Y(N112) );
  MXI4X1 U4402 ( .A(\block[0][1][30] ), .B(\block[1][1][30] ), .C(
        \block[2][1][30] ), .D(\block[3][1][30] ), .S0(n3616), .S1(n3645), .Y(
        n3470) );
  MXI4X1 U4403 ( .A(\block[4][1][30] ), .B(\block[5][1][30] ), .C(
        \block[6][1][30] ), .D(\block[7][1][30] ), .S0(n3608), .S1(n3645), .Y(
        n3471) );
  MXI2X1 U4404 ( .A(n3468), .B(n3469), .S0(n3662), .Y(N111) );
  MXI4X1 U4405 ( .A(\block[0][1][31] ), .B(\block[1][1][31] ), .C(
        \block[2][1][31] ), .D(\block[3][1][31] ), .S0(n3611), .S1(n3645), .Y(
        n3468) );
  MXI4X1 U4406 ( .A(\block[4][1][31] ), .B(\block[5][1][31] ), .C(
        \block[6][1][31] ), .D(\block[7][1][31] ), .S0(n3611), .S1(n3645), .Y(
        n3469) );
  OAI22XL U4407 ( .A0(n4148), .A1(n3858), .B0(n3868), .B1(n1122), .Y(n3169) );
  OAI22XL U4408 ( .A0(n4147), .A1(n3858), .B0(n3868), .B1(n1123), .Y(n3168) );
  OAI22XL U4409 ( .A0(n4146), .A1(n3858), .B0(n3868), .B1(n1124), .Y(n3167) );
  OAI22XL U4410 ( .A0(n4148), .A1(n3871), .B0(n3870), .B1(n1147), .Y(n3144) );
  OAI22XL U4411 ( .A0(n4147), .A1(n3871), .B0(n3880), .B1(n1148), .Y(n3143) );
  OAI22XL U4412 ( .A0(n4146), .A1(n3871), .B0(n3870), .B1(n1149), .Y(n3142) );
  OAI22XL U4413 ( .A0(n4148), .A1(n3884), .B0(n3894), .B1(n1172), .Y(n3119) );
  OAI22XL U4414 ( .A0(n4147), .A1(n3883), .B0(n3894), .B1(n1173), .Y(n3118) );
  OAI22XL U4415 ( .A0(n4146), .A1(n3883), .B0(n3894), .B1(n1174), .Y(n3117) );
  OAI22XL U4416 ( .A0(n4148), .A1(n3898), .B0(n3907), .B1(n1197), .Y(n3094) );
  OAI22XL U4417 ( .A0(n4147), .A1(n3897), .B0(n3907), .B1(n1198), .Y(n3093) );
  OAI22XL U4418 ( .A0(n4146), .A1(n3897), .B0(n3907), .B1(n1199), .Y(n3092) );
  OAI22XL U4419 ( .A0(n4148), .A1(n3911), .B0(n3920), .B1(n1222), .Y(n3069) );
  OAI22XL U4420 ( .A0(n4147), .A1(n3910), .B0(n3920), .B1(n1223), .Y(n3068) );
  OAI22XL U4421 ( .A0(n4146), .A1(n3910), .B0(n3920), .B1(n1224), .Y(n3067) );
  OAI22XL U4422 ( .A0(n4148), .A1(n3924), .B0(n3933), .B1(n1247), .Y(n3044) );
  OAI22XL U4423 ( .A0(n4147), .A1(n3923), .B0(n3933), .B1(n1248), .Y(n3043) );
  OAI22XL U4424 ( .A0(n4146), .A1(n3923), .B0(n3933), .B1(n1249), .Y(n3042) );
  OAI22XL U4425 ( .A0(n4148), .A1(n3937), .B0(n3946), .B1(n1272), .Y(n3019) );
  OAI22XL U4426 ( .A0(n4147), .A1(n3936), .B0(n3946), .B1(n1273), .Y(n3018) );
  OAI22XL U4427 ( .A0(n4146), .A1(n3936), .B0(n3946), .B1(n1274), .Y(n3017) );
  OAI22XL U4428 ( .A0(n4148), .A1(n3950), .B0(n3959), .B1(n1297), .Y(n2994) );
  OAI22XL U4429 ( .A0(n4147), .A1(n3949), .B0(n3959), .B1(n1298), .Y(n2993) );
  OAI22XL U4430 ( .A0(n4146), .A1(n3949), .B0(n3959), .B1(n1299), .Y(n2992) );
  OAI22XL U4431 ( .A0(n4145), .A1(n3858), .B0(n3868), .B1(n1125), .Y(n3166) );
  OAI22XL U4432 ( .A0(n4144), .A1(n3858), .B0(n3868), .B1(n1126), .Y(n3165) );
  OAI22XL U4433 ( .A0(n4143), .A1(n3858), .B0(n3868), .B1(n1127), .Y(n3164) );
  OAI22XL U4434 ( .A0(n4142), .A1(n3858), .B0(n3868), .B1(n1128), .Y(n3163) );
  OAI22XL U4435 ( .A0(n4141), .A1(n3858), .B0(n3867), .B1(n1129), .Y(n3162) );
  OAI22XL U4436 ( .A0(n4140), .A1(n3858), .B0(n3867), .B1(n1130), .Y(n3161) );
  OAI22XL U4437 ( .A0(n4139), .A1(n3858), .B0(n3868), .B1(n1131), .Y(n3160) );
  OAI22XL U4438 ( .A0(n4138), .A1(n3858), .B0(n3866), .B1(n1132), .Y(n3159) );
  OAI22XL U4439 ( .A0(n4137), .A1(n3858), .B0(n3868), .B1(n1133), .Y(n3158) );
  OAI22XL U4440 ( .A0(n4136), .A1(n3859), .B0(n3868), .B1(n1134), .Y(n3157) );
  OAI22XL U4441 ( .A0(n4135), .A1(n3859), .B0(n3866), .B1(n1135), .Y(n3156) );
  OAI22XL U4442 ( .A0(n4134), .A1(n3859), .B0(n3866), .B1(n1136), .Y(n3155) );
  OAI22XL U4443 ( .A0(n4133), .A1(n3859), .B0(n3866), .B1(n1137), .Y(n3154) );
  OAI22XL U4444 ( .A0(n4132), .A1(n3859), .B0(n3866), .B1(n1138), .Y(n3153) );
  OAI22XL U4445 ( .A0(n4131), .A1(n3859), .B0(n3866), .B1(n1139), .Y(n3152) );
  OAI22XL U4446 ( .A0(n4130), .A1(n3859), .B0(n3866), .B1(n1140), .Y(n3151) );
  OAI22XL U4447 ( .A0(n4129), .A1(n3859), .B0(n3868), .B1(n1141), .Y(n3150) );
  OAI22XL U4448 ( .A0(n4128), .A1(n3859), .B0(n3866), .B1(n1142), .Y(n3149) );
  OAI22XL U4449 ( .A0(n4127), .A1(n3859), .B0(n3866), .B1(n1143), .Y(n3148) );
  OAI22XL U4450 ( .A0(n4126), .A1(n3859), .B0(n3866), .B1(n1144), .Y(n3147) );
  OAI22XL U4451 ( .A0(n4125), .A1(n3859), .B0(n3868), .B1(n1145), .Y(n3146) );
  OAI22XL U4452 ( .A0(n4124), .A1(n3860), .B0(n3868), .B1(n1146), .Y(n3145) );
  OAI22XL U4453 ( .A0(n4145), .A1(n3871), .B0(n3870), .B1(n1150), .Y(n3141) );
  OAI22XL U4454 ( .A0(n4144), .A1(n3871), .B0(n3870), .B1(n1151), .Y(n3140) );
  OAI22XL U4455 ( .A0(n4143), .A1(n3871), .B0(n3880), .B1(n1152), .Y(n3139) );
  OAI22XL U4456 ( .A0(n4142), .A1(n3871), .B0(n3870), .B1(n1153), .Y(n3138) );
  OAI22XL U4457 ( .A0(n4141), .A1(n3871), .B0(n3881), .B1(n1154), .Y(n3137) );
  OAI22XL U4458 ( .A0(n4140), .A1(n3871), .B0(n3881), .B1(n1155), .Y(n3136) );
  OAI22XL U4459 ( .A0(n4139), .A1(n3871), .B0(n284), .B1(n1156), .Y(n3135) );
  OAI22XL U4460 ( .A0(n4138), .A1(n3871), .B0(n284), .B1(n1157), .Y(n3134) );
  OAI22XL U4461 ( .A0(n4137), .A1(n3871), .B0(n3870), .B1(n1158), .Y(n3133) );
  OAI22XL U4462 ( .A0(n4136), .A1(n3874), .B0(n3870), .B1(n1159), .Y(n3132) );
  OAI22XL U4463 ( .A0(n4135), .A1(n3873), .B0(n3880), .B1(n1160), .Y(n3131) );
  OAI22XL U4464 ( .A0(n4134), .A1(n3871), .B0(n3880), .B1(n1161), .Y(n3130) );
  OAI22XL U4465 ( .A0(n4133), .A1(n3874), .B0(n3880), .B1(n1162), .Y(n3129) );
  OAI22XL U4466 ( .A0(n4132), .A1(n3873), .B0(n3880), .B1(n1163), .Y(n3128) );
  OAI22XL U4467 ( .A0(n4131), .A1(n3871), .B0(n3880), .B1(n1164), .Y(n3127) );
  OAI22XL U4468 ( .A0(n4130), .A1(n3876), .B0(n3880), .B1(n1165), .Y(n3126) );
  OAI22XL U4469 ( .A0(n4129), .A1(n3874), .B0(n3880), .B1(n1166), .Y(n3125) );
  OAI22XL U4470 ( .A0(n4128), .A1(n3873), .B0(n3880), .B1(n1167), .Y(n3124) );
  OAI22XL U4471 ( .A0(n4127), .A1(n3873), .B0(n3870), .B1(n1168), .Y(n3123) );
  OAI22XL U4472 ( .A0(n4126), .A1(n3878), .B0(n3880), .B1(n1169), .Y(n3122) );
  OAI22XL U4473 ( .A0(n4125), .A1(n3874), .B0(n284), .B1(n1170), .Y(n3121) );
  OAI22XL U4474 ( .A0(n4124), .A1(n3872), .B0(n3880), .B1(n1171), .Y(n3120) );
  OAI22XL U4475 ( .A0(n4145), .A1(n3883), .B0(n3894), .B1(n1175), .Y(n3116) );
  OAI22XL U4476 ( .A0(n4144), .A1(n3891), .B0(n3894), .B1(n1176), .Y(n3115) );
  OAI22XL U4477 ( .A0(n4143), .A1(n3883), .B0(n3894), .B1(n1177), .Y(n3114) );
  OAI22XL U4478 ( .A0(n4142), .A1(n3883), .B0(n3894), .B1(n1178), .Y(n3113) );
  OAI22XL U4479 ( .A0(n4141), .A1(n3891), .B0(n3893), .B1(n1179), .Y(n3112) );
  OAI22XL U4480 ( .A0(n4140), .A1(n3883), .B0(n3893), .B1(n1180), .Y(n3111) );
  OAI22XL U4481 ( .A0(n4139), .A1(n3883), .B0(n3894), .B1(n1181), .Y(n3110) );
  OAI22XL U4482 ( .A0(n4138), .A1(n3891), .B0(n3894), .B1(n1182), .Y(n3109) );
  OAI22XL U4483 ( .A0(n4137), .A1(n3883), .B0(n3892), .B1(n1183), .Y(n3108) );
  OAI22XL U4484 ( .A0(n4136), .A1(n3883), .B0(n3892), .B1(n1184), .Y(n3107) );
  OAI22XL U4485 ( .A0(n4135), .A1(n3883), .B0(n3892), .B1(n1185), .Y(n3106) );
  OAI22XL U4486 ( .A0(n4134), .A1(n3883), .B0(n3892), .B1(n1186), .Y(n3105) );
  OAI22XL U4487 ( .A0(n4133), .A1(n3883), .B0(n3894), .B1(n1187), .Y(n3104) );
  OAI22XL U4488 ( .A0(n4132), .A1(n3883), .B0(n3894), .B1(n1188), .Y(n3103) );
  OAI22XL U4489 ( .A0(n4131), .A1(n3883), .B0(n3894), .B1(n1189), .Y(n3102) );
  OAI22XL U4490 ( .A0(n4130), .A1(n3883), .B0(n3892), .B1(n1190), .Y(n3101) );
  OAI22XL U4491 ( .A0(n4129), .A1(n3883), .B0(n3892), .B1(n1191), .Y(n3100) );
  OAI22XL U4492 ( .A0(n4128), .A1(n3883), .B0(n3892), .B1(n1192), .Y(n3099) );
  OAI22XL U4493 ( .A0(n4127), .A1(n3891), .B0(n3894), .B1(n1193), .Y(n3098) );
  OAI22XL U4494 ( .A0(n4126), .A1(n3883), .B0(n3894), .B1(n1194), .Y(n3097) );
  OAI22XL U4495 ( .A0(n4125), .A1(n3883), .B0(n3892), .B1(n1195), .Y(n3096) );
  OAI22XL U4496 ( .A0(n4124), .A1(n3891), .B0(n3892), .B1(n1196), .Y(n3095) );
  OAI22XL U4497 ( .A0(n4145), .A1(n3897), .B0(n3907), .B1(n1200), .Y(n3091) );
  OAI22XL U4498 ( .A0(n4144), .A1(n3897), .B0(n3907), .B1(n1201), .Y(n3090) );
  OAI22XL U4499 ( .A0(n4143), .A1(n3897), .B0(n3907), .B1(n1202), .Y(n3089) );
  OAI22XL U4500 ( .A0(n4142), .A1(n3897), .B0(n3907), .B1(n1203), .Y(n3088) );
  OAI22XL U4501 ( .A0(n4141), .A1(n3897), .B0(n3906), .B1(n1204), .Y(n3087) );
  OAI22XL U4502 ( .A0(n4140), .A1(n3897), .B0(n3906), .B1(n1205), .Y(n3086) );
  OAI22XL U4503 ( .A0(n4139), .A1(n3897), .B0(n3907), .B1(n1206), .Y(n3085) );
  OAI22XL U4504 ( .A0(n4138), .A1(n3897), .B0(n3905), .B1(n1207), .Y(n3084) );
  OAI22XL U4505 ( .A0(n4137), .A1(n3897), .B0(n3907), .B1(n1208), .Y(n3083) );
  OAI22XL U4506 ( .A0(n4136), .A1(n3897), .B0(n3907), .B1(n1209), .Y(n3082) );
  OAI22XL U4507 ( .A0(n4135), .A1(n3902), .B0(n3905), .B1(n1210), .Y(n3081) );
  OAI22XL U4508 ( .A0(n4134), .A1(n3901), .B0(n3905), .B1(n1211), .Y(n3080) );
  OAI22XL U4509 ( .A0(n4133), .A1(n3900), .B0(n3905), .B1(n1212), .Y(n3079) );
  OAI22XL U4510 ( .A0(n4132), .A1(n3902), .B0(n3905), .B1(n1213), .Y(n3078) );
  OAI22XL U4511 ( .A0(n4131), .A1(n3901), .B0(n3905), .B1(n1214), .Y(n3077) );
  OAI22XL U4512 ( .A0(n4130), .A1(n3900), .B0(n3905), .B1(n1215), .Y(n3076) );
  OAI22XL U4513 ( .A0(n4129), .A1(n3902), .B0(n3905), .B1(n1216), .Y(n3075) );
  OAI22XL U4514 ( .A0(n4128), .A1(n3901), .B0(n3905), .B1(n1217), .Y(n3074) );
  OAI22XL U4515 ( .A0(n4127), .A1(n3898), .B0(n3905), .B1(n1218), .Y(n3073) );
  OAI22XL U4516 ( .A0(n4126), .A1(n3899), .B0(n3907), .B1(n1219), .Y(n3072) );
  OAI22XL U4517 ( .A0(n4125), .A1(n3904), .B0(n3907), .B1(n1220), .Y(n3071) );
  OAI22XL U4518 ( .A0(n4124), .A1(n3900), .B0(n3907), .B1(n1221), .Y(n3070) );
  OAI22XL U4519 ( .A0(n4145), .A1(n3910), .B0(n3920), .B1(n1225), .Y(n3066) );
  OAI22XL U4520 ( .A0(n4144), .A1(n3910), .B0(n3920), .B1(n1226), .Y(n3065) );
  OAI22XL U4521 ( .A0(n4143), .A1(n3910), .B0(n3920), .B1(n1227), .Y(n3064) );
  OAI22XL U4522 ( .A0(n4142), .A1(n3910), .B0(n3920), .B1(n1228), .Y(n3063) );
  OAI22XL U4523 ( .A0(n4141), .A1(n3910), .B0(n3919), .B1(n1229), .Y(n3062) );
  OAI22XL U4524 ( .A0(n4140), .A1(n3910), .B0(n3919), .B1(n1230), .Y(n3061) );
  OAI22XL U4525 ( .A0(n4139), .A1(n3910), .B0(n3918), .B1(n1231), .Y(n3060) );
  OAI22XL U4526 ( .A0(n4138), .A1(n3910), .B0(n3918), .B1(n1232), .Y(n3059) );
  OAI22XL U4527 ( .A0(n4137), .A1(n3910), .B0(n3920), .B1(n1233), .Y(n3058) );
  OAI22XL U4528 ( .A0(n4136), .A1(n3910), .B0(n3920), .B1(n1234), .Y(n3057) );
  OAI22XL U4529 ( .A0(n4135), .A1(n3913), .B0(n3918), .B1(n1235), .Y(n3056) );
  OAI22XL U4530 ( .A0(n4134), .A1(n3914), .B0(n3918), .B1(n1236), .Y(n3055) );
  OAI22XL U4531 ( .A0(n4133), .A1(n3915), .B0(n3918), .B1(n1237), .Y(n3054) );
  OAI22XL U4532 ( .A0(n4132), .A1(n3913), .B0(n3918), .B1(n1238), .Y(n3053) );
  OAI22XL U4533 ( .A0(n4131), .A1(n3914), .B0(n3918), .B1(n1239), .Y(n3052) );
  OAI22XL U4534 ( .A0(n4130), .A1(n3915), .B0(n3918), .B1(n1240), .Y(n3051) );
  OAI22XL U4535 ( .A0(n4129), .A1(n3913), .B0(n3918), .B1(n1241), .Y(n3050) );
  OAI22XL U4536 ( .A0(n4128), .A1(n3912), .B0(n3920), .B1(n1242), .Y(n3049) );
  OAI22XL U4537 ( .A0(n4127), .A1(n3911), .B0(n3918), .B1(n1243), .Y(n3048) );
  OAI22XL U4538 ( .A0(n4126), .A1(n3917), .B0(n3920), .B1(n1244), .Y(n3047) );
  OAI22XL U4539 ( .A0(n4125), .A1(n3914), .B0(n3920), .B1(n1245), .Y(n3046) );
  OAI22XL U4540 ( .A0(n4124), .A1(n3915), .B0(n3920), .B1(n1246), .Y(n3045) );
  OAI22XL U4541 ( .A0(n4145), .A1(n3923), .B0(n3933), .B1(n1250), .Y(n3041) );
  OAI22XL U4542 ( .A0(n4144), .A1(n3923), .B0(n3933), .B1(n1251), .Y(n3040) );
  OAI22XL U4543 ( .A0(n4143), .A1(n3923), .B0(n3933), .B1(n1252), .Y(n3039) );
  OAI22XL U4544 ( .A0(n4142), .A1(n3923), .B0(n3933), .B1(n1253), .Y(n3038) );
  OAI22XL U4545 ( .A0(n4141), .A1(n3923), .B0(n3932), .B1(n1254), .Y(n3037) );
  OAI22XL U4546 ( .A0(n4140), .A1(n3923), .B0(n3932), .B1(n1255), .Y(n3036) );
  OAI22XL U4547 ( .A0(n4139), .A1(n3923), .B0(n3931), .B1(n1256), .Y(n3035) );
  OAI22XL U4548 ( .A0(n4138), .A1(n3923), .B0(n3931), .B1(n1257), .Y(n3034) );
  OAI22XL U4549 ( .A0(n4137), .A1(n3923), .B0(n3933), .B1(n1258), .Y(n3033) );
  OAI22XL U4550 ( .A0(n4136), .A1(n3923), .B0(n3933), .B1(n1259), .Y(n3032) );
  OAI22XL U4551 ( .A0(n4135), .A1(n3926), .B0(n3931), .B1(n1260), .Y(n3031) );
  OAI22XL U4552 ( .A0(n4134), .A1(n3927), .B0(n3931), .B1(n1261), .Y(n3030) );
  OAI22XL U4553 ( .A0(n4133), .A1(n3928), .B0(n3931), .B1(n1262), .Y(n3029) );
  OAI22XL U4554 ( .A0(n4132), .A1(n3926), .B0(n3931), .B1(n1263), .Y(n3028) );
  OAI22XL U4555 ( .A0(n4131), .A1(n3927), .B0(n3931), .B1(n1264), .Y(n3027) );
  OAI22XL U4556 ( .A0(n4130), .A1(n3928), .B0(n3931), .B1(n1265), .Y(n3026) );
  OAI22XL U4557 ( .A0(n4129), .A1(n3926), .B0(n3931), .B1(n1266), .Y(n3025) );
  OAI22XL U4558 ( .A0(n4128), .A1(n3925), .B0(n3933), .B1(n1267), .Y(n3024) );
  OAI22XL U4559 ( .A0(n4127), .A1(n3924), .B0(n3931), .B1(n1268), .Y(n3023) );
  OAI22XL U4560 ( .A0(n4126), .A1(n3930), .B0(n3933), .B1(n1269), .Y(n3022) );
  OAI22XL U4561 ( .A0(n4125), .A1(n3927), .B0(n3933), .B1(n1270), .Y(n3021) );
  OAI22XL U4562 ( .A0(n4124), .A1(n3928), .B0(n3933), .B1(n1271), .Y(n3020) );
  OAI22XL U4563 ( .A0(n4145), .A1(n3936), .B0(n3946), .B1(n1275), .Y(n3016) );
  OAI22XL U4564 ( .A0(n4144), .A1(n3936), .B0(n3946), .B1(n1276), .Y(n3015) );
  OAI22XL U4565 ( .A0(n4143), .A1(n3936), .B0(n3946), .B1(n1277), .Y(n3014) );
  OAI22XL U4566 ( .A0(n4142), .A1(n3936), .B0(n3946), .B1(n1278), .Y(n3013) );
  OAI22XL U4567 ( .A0(n4141), .A1(n3936), .B0(n3945), .B1(n1279), .Y(n3012) );
  OAI22XL U4568 ( .A0(n4140), .A1(n3936), .B0(n3945), .B1(n1280), .Y(n3011) );
  OAI22XL U4569 ( .A0(n4139), .A1(n3936), .B0(n3944), .B1(n1281), .Y(n3010) );
  OAI22XL U4570 ( .A0(n4138), .A1(n3936), .B0(n3944), .B1(n1282), .Y(n3009) );
  OAI22XL U4571 ( .A0(n4137), .A1(n3936), .B0(n3946), .B1(n1283), .Y(n3008) );
  OAI22XL U4572 ( .A0(n4136), .A1(n3936), .B0(n3946), .B1(n1284), .Y(n3007) );
  OAI22XL U4573 ( .A0(n4135), .A1(n3939), .B0(n3944), .B1(n1285), .Y(n3006) );
  OAI22XL U4574 ( .A0(n4134), .A1(n3940), .B0(n3944), .B1(n1286), .Y(n3005) );
  OAI22XL U4575 ( .A0(n4133), .A1(n3941), .B0(n3944), .B1(n1287), .Y(n3004) );
  OAI22XL U4576 ( .A0(n4132), .A1(n3939), .B0(n3944), .B1(n1288), .Y(n3003) );
  OAI22XL U4577 ( .A0(n4131), .A1(n3940), .B0(n3944), .B1(n1289), .Y(n3002) );
  OAI22XL U4578 ( .A0(n4130), .A1(n3941), .B0(n3944), .B1(n1290), .Y(n3001) );
  OAI22XL U4579 ( .A0(n4129), .A1(n3939), .B0(n3944), .B1(n1291), .Y(n3000) );
  OAI22XL U4580 ( .A0(n4128), .A1(n3938), .B0(n3946), .B1(n1292), .Y(n2999) );
  OAI22XL U4581 ( .A0(n4127), .A1(n3937), .B0(n3944), .B1(n1293), .Y(n2998) );
  OAI22XL U4582 ( .A0(n4126), .A1(n3943), .B0(n3946), .B1(n1294), .Y(n2997) );
  OAI22XL U4583 ( .A0(n4125), .A1(n3940), .B0(n3946), .B1(n1295), .Y(n2996) );
  OAI22XL U4584 ( .A0(n4124), .A1(n3941), .B0(n3946), .B1(n1296), .Y(n2995) );
  OAI22XL U4585 ( .A0(n4145), .A1(n3949), .B0(n3959), .B1(n1300), .Y(n2991) );
  OAI22XL U4586 ( .A0(n4144), .A1(n3949), .B0(n3959), .B1(n1301), .Y(n2990) );
  OAI22XL U4587 ( .A0(n4143), .A1(n3949), .B0(n3959), .B1(n1302), .Y(n2989) );
  OAI22XL U4588 ( .A0(n4142), .A1(n3949), .B0(n3959), .B1(n1303), .Y(n2988) );
  OAI22XL U4589 ( .A0(n4141), .A1(n3949), .B0(n3958), .B1(n1304), .Y(n2987) );
  OAI22XL U4590 ( .A0(n4140), .A1(n3949), .B0(n3958), .B1(n1305), .Y(n2986) );
  OAI22XL U4591 ( .A0(n4139), .A1(n3949), .B0(n3957), .B1(n1306), .Y(n2985) );
  OAI22XL U4592 ( .A0(n4138), .A1(n3949), .B0(n3957), .B1(n1307), .Y(n2984) );
  OAI22XL U4593 ( .A0(n4137), .A1(n3949), .B0(n3959), .B1(n1308), .Y(n2983) );
  OAI22XL U4594 ( .A0(n4136), .A1(n3949), .B0(n3959), .B1(n1309), .Y(n2982) );
  OAI22XL U4595 ( .A0(n4135), .A1(n3953), .B0(n3957), .B1(n1310), .Y(n2981) );
  OAI22XL U4596 ( .A0(n4134), .A1(n3952), .B0(n3957), .B1(n1311), .Y(n2980) );
  OAI22XL U4597 ( .A0(n4133), .A1(n3954), .B0(n3957), .B1(n1312), .Y(n2979) );
  OAI22XL U4598 ( .A0(n4132), .A1(n3953), .B0(n3957), .B1(n1313), .Y(n2978) );
  OAI22XL U4599 ( .A0(n4131), .A1(n3952), .B0(n3957), .B1(n1314), .Y(n2977) );
  OAI22XL U4600 ( .A0(n4130), .A1(n3954), .B0(n3957), .B1(n1315), .Y(n2976) );
  OAI22XL U4601 ( .A0(n4129), .A1(n3953), .B0(n3957), .B1(n1316), .Y(n2975) );
  OAI22XL U4602 ( .A0(n4128), .A1(n3951), .B0(n3959), .B1(n1317), .Y(n2974) );
  OAI22XL U4603 ( .A0(n4127), .A1(n3950), .B0(n3957), .B1(n1318), .Y(n2973) );
  OAI22XL U4604 ( .A0(n4126), .A1(n3956), .B0(n3959), .B1(n1319), .Y(n2972) );
  OAI22XL U4605 ( .A0(n4125), .A1(n3952), .B0(n3959), .B1(n1320), .Y(n2971) );
  OAI22XL U4606 ( .A0(n4124), .A1(n3954), .B0(n3959), .B1(n1321), .Y(n2970) );
  NAND3X1 U4607 ( .A(n3807), .B(n303), .C(proc_read), .Y(n200) );
  NAND2X1 U4608 ( .A(n1703), .B(n3860), .Y(n1704) );
  NAND2X1 U4609 ( .A(n1702), .B(n3872), .Y(n1705) );
  NAND2X1 U4610 ( .A(n1700), .B(n3898), .Y(n1707) );
  NAND2X1 U4611 ( .A(n1699), .B(n3911), .Y(n1708) );
  NAND2X1 U4612 ( .A(n1698), .B(n3924), .Y(n1709) );
  NAND2X1 U4613 ( .A(n1697), .B(n3937), .Y(n1710) );
  NAND2X1 U4614 ( .A(n1696), .B(n3950), .Y(n1711) );
  NAND2X1 U4615 ( .A(n1701), .B(n3884), .Y(n1706) );
  AO22X1 U4616 ( .A0(n4000), .A1(next_proc_wdata[0]), .B0(n4002), .B1(
        proc_wdata[0]), .Y(n2812) );
  AO22X1 U4617 ( .A0(n4000), .A1(next_proc_wdata[1]), .B0(n4002), .B1(
        proc_wdata[1]), .Y(n2811) );
  AO22X1 U4618 ( .A0(n4000), .A1(next_proc_wdata[2]), .B0(n4002), .B1(
        proc_wdata[2]), .Y(n2810) );
  AO22X1 U4619 ( .A0(n4000), .A1(next_proc_wdata[3]), .B0(n4002), .B1(
        proc_wdata[3]), .Y(n2809) );
  AO22X1 U4620 ( .A0(n4000), .A1(next_proc_wdata[4]), .B0(n4002), .B1(
        proc_wdata[4]), .Y(n2808) );
  AO22X1 U4621 ( .A0(n4000), .A1(next_proc_wdata[5]), .B0(n4002), .B1(
        proc_wdata[5]), .Y(n2807) );
  AO22X1 U4622 ( .A0(n4000), .A1(next_proc_wdata[6]), .B0(n3281), .B1(
        proc_wdata[6]), .Y(n2806) );
  AO22X1 U4623 ( .A0(n4000), .A1(next_proc_wdata[7]), .B0(n3281), .B1(
        proc_wdata[7]), .Y(n2805) );
  AO22X1 U4624 ( .A0(n4000), .A1(next_proc_wdata[8]), .B0(n3281), .B1(
        proc_wdata[8]), .Y(n2804) );
  AO22X1 U4625 ( .A0(n4000), .A1(next_proc_wdata[9]), .B0(n3281), .B1(
        proc_wdata[9]), .Y(n2803) );
  AO22X1 U4626 ( .A0(n4000), .A1(next_proc_wdata[10]), .B0(n3281), .B1(
        proc_wdata[10]), .Y(n2802) );
  AO22X1 U4627 ( .A0(n4000), .A1(next_proc_wdata[11]), .B0(n3281), .B1(
        proc_wdata[11]), .Y(n2801) );
  AO22X1 U4628 ( .A0(n4000), .A1(next_proc_wdata[12]), .B0(n4002), .B1(
        proc_wdata[12]), .Y(n2800) );
  AO22X1 U4629 ( .A0(n4000), .A1(next_proc_wdata[13]), .B0(n4002), .B1(
        proc_wdata[13]), .Y(n2799) );
  AO22X1 U4630 ( .A0(n4001), .A1(next_proc_wdata[14]), .B0(n4002), .B1(
        proc_wdata[14]), .Y(n2798) );
  AO22X1 U4631 ( .A0(n4001), .A1(next_proc_wdata[15]), .B0(n4002), .B1(
        proc_wdata[15]), .Y(n2797) );
  AO22X1 U4632 ( .A0(n4001), .A1(next_proc_wdata[16]), .B0(n4002), .B1(
        proc_wdata[16]), .Y(n2796) );
  AO22X1 U4633 ( .A0(n4001), .A1(next_proc_wdata[17]), .B0(n4002), .B1(
        proc_wdata[17]), .Y(n2795) );
  AO22X1 U4634 ( .A0(n4001), .A1(next_proc_wdata[18]), .B0(n4002), .B1(
        proc_wdata[18]), .Y(n2794) );
  AO22X1 U4635 ( .A0(n4001), .A1(next_proc_wdata[19]), .B0(n4002), .B1(
        proc_wdata[19]), .Y(n2793) );
  AO22X1 U4636 ( .A0(n4001), .A1(next_proc_wdata[20]), .B0(n3281), .B1(
        proc_wdata[20]), .Y(n2792) );
  AO22X1 U4637 ( .A0(n4001), .A1(next_proc_wdata[21]), .B0(n4002), .B1(
        proc_wdata[21]), .Y(n2791) );
  AO22X1 U4638 ( .A0(n4001), .A1(next_proc_wdata[22]), .B0(n3281), .B1(
        proc_wdata[22]), .Y(n2790) );
  AO22X1 U4639 ( .A0(n4001), .A1(next_proc_wdata[23]), .B0(n4002), .B1(
        proc_wdata[23]), .Y(n2789) );
  AO22X1 U4640 ( .A0(n4001), .A1(next_proc_wdata[24]), .B0(n3281), .B1(
        proc_wdata[24]), .Y(n2788) );
  AO22X1 U4641 ( .A0(n4001), .A1(next_proc_wdata[25]), .B0(n4002), .B1(
        proc_wdata[25]), .Y(n2787) );
  AO22X1 U4642 ( .A0(n4001), .A1(next_proc_wdata[26]), .B0(n3281), .B1(
        proc_wdata[26]), .Y(n2786) );
  AO22X1 U4643 ( .A0(n4001), .A1(next_proc_wdata[27]), .B0(n4002), .B1(
        proc_wdata[27]), .Y(n2785) );
  AO22X1 U4644 ( .A0(n4001), .A1(next_proc_wdata[28]), .B0(n4002), .B1(
        proc_wdata[28]), .Y(n2784) );
  AO22X1 U4645 ( .A0(n4001), .A1(next_proc_wdata[29]), .B0(n3281), .B1(
        proc_wdata[29]), .Y(n2783) );
  AO22X1 U4646 ( .A0(n4001), .A1(next_proc_wdata[30]), .B0(n3281), .B1(
        proc_wdata[30]), .Y(n2782) );
  AO22X1 U4647 ( .A0(n4001), .A1(next_proc_wdata[31]), .B0(n4002), .B1(
        proc_wdata[31]), .Y(n2781) );
  INVX3 U4648 ( .A(mem_rdata[57]), .Y(n4245) );
  INVX3 U4649 ( .A(mem_rdata[58]), .Y(n4244) );
  INVX3 U4650 ( .A(mem_rdata[59]), .Y(n4243) );
  INVX3 U4651 ( .A(mem_rdata[60]), .Y(n4242) );
  INVX3 U4652 ( .A(mem_rdata[61]), .Y(n4241) );
  INVX3 U4653 ( .A(mem_rdata[62]), .Y(n4240) );
  INVX3 U4654 ( .A(mem_rdata[63]), .Y(n4239) );
  INVX3 U4655 ( .A(mem_rdata[64]), .Y(n4238) );
  INVX3 U4656 ( .A(mem_rdata[65]), .Y(n4237) );
  INVX3 U4657 ( .A(mem_rdata[66]), .Y(n4236) );
  INVX3 U4658 ( .A(mem_rdata[67]), .Y(n4235) );
  INVX3 U4659 ( .A(mem_rdata[68]), .Y(n4234) );
  INVX3 U4660 ( .A(mem_rdata[69]), .Y(n4233) );
  INVX3 U4661 ( .A(mem_rdata[70]), .Y(n4232) );
  INVX3 U4662 ( .A(mem_rdata[71]), .Y(n4231) );
  INVX3 U4663 ( .A(mem_rdata[72]), .Y(n4230) );
  INVX3 U4664 ( .A(mem_rdata[73]), .Y(n4229) );
  INVX3 U4665 ( .A(mem_rdata[74]), .Y(n4228) );
  INVX3 U4666 ( .A(mem_rdata[75]), .Y(n4227) );
  INVX3 U4667 ( .A(mem_rdata[76]), .Y(n4226) );
  INVX3 U4668 ( .A(mem_rdata[77]), .Y(n4225) );
  INVX3 U4669 ( .A(mem_rdata[78]), .Y(n4224) );
  INVX3 U4670 ( .A(mem_rdata[79]), .Y(n4223) );
  INVX3 U4671 ( .A(mem_rdata[80]), .Y(n4222) );
  INVX3 U4672 ( .A(mem_rdata[81]), .Y(n4221) );
  INVX3 U4673 ( .A(mem_rdata[82]), .Y(n4220) );
  INVX3 U4674 ( .A(mem_rdata[83]), .Y(n4219) );
  INVX3 U4675 ( .A(mem_rdata[84]), .Y(n4218) );
  INVX3 U4676 ( .A(mem_rdata[85]), .Y(n4217) );
  INVX3 U4677 ( .A(mem_rdata[86]), .Y(n4216) );
  INVX3 U4678 ( .A(mem_rdata[87]), .Y(n4215) );
  INVX3 U4679 ( .A(mem_rdata[88]), .Y(n4214) );
  INVX3 U4680 ( .A(mem_rdata[89]), .Y(n4213) );
  INVX3 U4681 ( .A(mem_rdata[90]), .Y(n4212) );
  INVX3 U4682 ( .A(mem_rdata[91]), .Y(n4211) );
  INVX3 U4683 ( .A(mem_rdata[92]), .Y(n4210) );
  INVX3 U4684 ( .A(mem_rdata[93]), .Y(n4209) );
  INVX3 U4685 ( .A(mem_rdata[94]), .Y(n4208) );
  INVX3 U4686 ( .A(mem_rdata[95]), .Y(n4207) );
  INVX3 U4687 ( .A(mem_rdata[96]), .Y(n4206) );
  INVX3 U4688 ( .A(mem_rdata[97]), .Y(n4205) );
  INVX3 U4689 ( .A(mem_rdata[98]), .Y(n4204) );
  INVX3 U4690 ( .A(mem_rdata[99]), .Y(n4203) );
  INVX3 U4691 ( .A(mem_rdata[100]), .Y(n4202) );
  INVX3 U4692 ( .A(mem_rdata[101]), .Y(n4201) );
  INVX3 U4693 ( .A(mem_rdata[102]), .Y(n4200) );
  INVX3 U4694 ( .A(mem_rdata[103]), .Y(n4199) );
  INVX3 U4695 ( .A(mem_rdata[104]), .Y(n4198) );
  INVX3 U4696 ( .A(mem_rdata[105]), .Y(n4197) );
  INVX3 U4697 ( .A(mem_rdata[106]), .Y(n4196) );
  INVX3 U4698 ( .A(mem_rdata[107]), .Y(n4195) );
  INVX3 U4699 ( .A(mem_rdata[108]), .Y(n4194) );
  INVX3 U4700 ( .A(mem_rdata[109]), .Y(n4193) );
  INVX3 U4701 ( .A(mem_rdata[110]), .Y(n4192) );
  INVX3 U4702 ( .A(mem_rdata[111]), .Y(n4191) );
  INVX3 U4703 ( .A(mem_rdata[112]), .Y(n4190) );
  INVX3 U4704 ( .A(mem_rdata[113]), .Y(n4189) );
  INVX3 U4705 ( .A(mem_rdata[114]), .Y(n4188) );
  INVX3 U4706 ( .A(mem_rdata[115]), .Y(n4187) );
  INVX3 U4707 ( .A(mem_rdata[116]), .Y(n4186) );
  INVX3 U4708 ( .A(mem_rdata[117]), .Y(n4185) );
  INVX3 U4709 ( .A(mem_rdata[118]), .Y(n4184) );
  INVX3 U4710 ( .A(mem_rdata[119]), .Y(n4183) );
  INVX3 U4711 ( .A(mem_rdata[120]), .Y(n4182) );
  INVX3 U4712 ( .A(mem_rdata[121]), .Y(n4181) );
  INVX3 U4713 ( .A(mem_rdata[122]), .Y(n4180) );
  INVX3 U4714 ( .A(mem_rdata[123]), .Y(n4179) );
  INVX3 U4715 ( .A(mem_rdata[124]), .Y(n4178) );
  INVX3 U4716 ( .A(mem_rdata[125]), .Y(n4177) );
  INVX3 U4717 ( .A(mem_rdata[126]), .Y(n4176) );
  INVX3 U4718 ( .A(mem_rdata[127]), .Y(n4175) );
  INVX3 U4719 ( .A(mem_rdata[32]), .Y(n4270) );
  INVX3 U4720 ( .A(mem_rdata[33]), .Y(n4269) );
  INVX3 U4721 ( .A(mem_rdata[34]), .Y(n4268) );
  INVX3 U4722 ( .A(mem_rdata[35]), .Y(n4267) );
  INVX3 U4723 ( .A(mem_rdata[36]), .Y(n4266) );
  INVX3 U4724 ( .A(mem_rdata[37]), .Y(n4265) );
  INVX3 U4725 ( .A(mem_rdata[38]), .Y(n4264) );
  INVX3 U4726 ( .A(mem_rdata[39]), .Y(n4263) );
  INVX3 U4727 ( .A(mem_rdata[40]), .Y(n4262) );
  INVX3 U4728 ( .A(mem_rdata[41]), .Y(n4261) );
  INVX3 U4729 ( .A(mem_rdata[42]), .Y(n4260) );
  INVX3 U4730 ( .A(mem_rdata[43]), .Y(n4259) );
  INVX3 U4731 ( .A(mem_rdata[44]), .Y(n4258) );
  INVX3 U4732 ( .A(mem_rdata[45]), .Y(n4257) );
  INVX3 U4733 ( .A(mem_rdata[46]), .Y(n4256) );
  INVX3 U4734 ( .A(mem_rdata[47]), .Y(n4255) );
  INVX3 U4735 ( .A(mem_rdata[48]), .Y(n4254) );
  INVX3 U4736 ( .A(mem_rdata[49]), .Y(n4253) );
  INVX3 U4737 ( .A(mem_rdata[50]), .Y(n4252) );
  INVX3 U4738 ( .A(mem_rdata[51]), .Y(n4251) );
  INVX3 U4739 ( .A(mem_rdata[52]), .Y(n4250) );
  INVX3 U4740 ( .A(mem_rdata[53]), .Y(n4249) );
  INVX3 U4741 ( .A(mem_rdata[54]), .Y(n4248) );
  INVX3 U4742 ( .A(mem_rdata[55]), .Y(n4247) );
  INVX3 U4743 ( .A(mem_rdata[56]), .Y(n4246) );
  INVX3 U4744 ( .A(mem_rdata[0]), .Y(n4302) );
  INVX3 U4745 ( .A(mem_rdata[1]), .Y(n4301) );
  INVX3 U4746 ( .A(mem_rdata[2]), .Y(n4300) );
  INVX3 U4747 ( .A(mem_rdata[3]), .Y(n4299) );
  INVX3 U4748 ( .A(mem_rdata[4]), .Y(n4298) );
  INVX3 U4749 ( .A(mem_rdata[5]), .Y(n4297) );
  INVX3 U4750 ( .A(mem_rdata[6]), .Y(n4296) );
  INVX3 U4751 ( .A(mem_rdata[7]), .Y(n4295) );
  INVX3 U4752 ( .A(mem_rdata[8]), .Y(n4294) );
  INVX3 U4753 ( .A(mem_rdata[9]), .Y(n4293) );
  INVX3 U4754 ( .A(mem_rdata[10]), .Y(n4292) );
  INVX3 U4755 ( .A(mem_rdata[11]), .Y(n4291) );
  INVX3 U4756 ( .A(mem_rdata[12]), .Y(n4290) );
  INVX3 U4757 ( .A(mem_rdata[13]), .Y(n4289) );
  INVX3 U4758 ( .A(mem_rdata[14]), .Y(n4288) );
  INVX3 U4759 ( .A(mem_rdata[15]), .Y(n4287) );
  INVX3 U4760 ( .A(mem_rdata[16]), .Y(n4286) );
  INVX3 U4761 ( .A(mem_rdata[17]), .Y(n4285) );
  INVX3 U4762 ( .A(mem_rdata[18]), .Y(n4284) );
  INVX3 U4763 ( .A(mem_rdata[19]), .Y(n4283) );
  INVX3 U4764 ( .A(mem_rdata[20]), .Y(n4282) );
  INVX3 U4765 ( .A(mem_rdata[21]), .Y(n4281) );
  INVX3 U4766 ( .A(mem_rdata[22]), .Y(n4280) );
  INVX3 U4767 ( .A(mem_rdata[23]), .Y(n4279) );
  INVX3 U4768 ( .A(mem_rdata[24]), .Y(n4278) );
  INVX3 U4769 ( .A(mem_rdata[25]), .Y(n4277) );
  INVX3 U4770 ( .A(mem_rdata[26]), .Y(n4276) );
  INVX3 U4771 ( .A(mem_rdata[27]), .Y(n4275) );
  INVX3 U4772 ( .A(mem_rdata[28]), .Y(n4274) );
  INVX3 U4773 ( .A(mem_rdata[29]), .Y(n4273) );
  INVX3 U4774 ( .A(mem_rdata[30]), .Y(n4272) );
  INVX3 U4775 ( .A(mem_rdata[31]), .Y(n4271) );
  NAND2X1 U4776 ( .A(state[0]), .B(state[1]), .Y(n302) );
  INVX3 U4777 ( .A(proc_addr[5]), .Y(n4148) );
  INVX3 U4778 ( .A(proc_addr[6]), .Y(n4147) );
  INVX3 U4779 ( .A(proc_addr[8]), .Y(n4145) );
  INVX3 U4780 ( .A(proc_addr[13]), .Y(n4140) );
  INVX3 U4781 ( .A(proc_addr[14]), .Y(n4139) );
  INVX3 U4782 ( .A(proc_addr[15]), .Y(n4138) );
  INVX3 U4783 ( .A(proc_addr[16]), .Y(n4137) );
  INVX3 U4784 ( .A(proc_addr[17]), .Y(n4136) );
  INVX3 U4785 ( .A(proc_addr[18]), .Y(n4135) );
  INVX3 U4786 ( .A(proc_addr[19]), .Y(n4134) );
  INVX3 U4787 ( .A(proc_addr[20]), .Y(n4133) );
  INVX3 U4788 ( .A(proc_addr[24]), .Y(n4129) );
  INVX3 U4789 ( .A(proc_addr[25]), .Y(n4128) );
endmodule

